
module CONT ( clk, reset, im_wen_n, cr_a, curr_time, fb_addr, photo_num, 
        curr_photo_addr, curr_photo_size, en_si, en_init_time, en_fb_addr, 
        en_photo_num, en_curr_photo_addr, en_curr_photo_size, en_so, si_sel, 
        init_time_mux_sel, sftr_n, so_mux_sel, expand_sel, \im_a[19]_BAR , 
        \im_a[18]_BAR , \im_a[17]_BAR , \im_a[16]_BAR , \im_a[15]_BAR , 
        \im_a[14]_BAR , \im_a[13]_BAR , \im_a[12]_BAR , \im_a[11]_BAR , 
        \im_a[10]_BAR , \im_a[9]_BAR , \im_a[8]_BAR , \im_a[7]_BAR , 
        \im_a[6]_BAR , \im_a[5]_BAR , \im_a[4]_BAR , \im_a[3]_BAR , 
        \im_a[2]_BAR , \im_a[1]_BAR , \im_a[0]_BAR  );
  output [8:0] cr_a;
  input [23:0] curr_time;
  input [19:0] fb_addr;
  input [1:0] photo_num;
  input [19:0] curr_photo_addr;
  input [1:0] curr_photo_size;
  output [1:0] sftr_n;
  output [1:0] so_mux_sel;
  output [3:0] expand_sel;
  input clk, reset;
  output im_wen_n, en_si, en_init_time, en_fb_addr, en_photo_num,
         en_curr_photo_addr, en_curr_photo_size, en_so, si_sel,
         init_time_mux_sel, \im_a[19]_BAR , \im_a[18]_BAR , \im_a[17]_BAR ,
         \im_a[16]_BAR , \im_a[15]_BAR , \im_a[14]_BAR , \im_a[13]_BAR ,
         \im_a[12]_BAR , \im_a[11]_BAR , \im_a[10]_BAR , \im_a[9]_BAR ,
         \im_a[8]_BAR , \im_a[7]_BAR , \im_a[6]_BAR , \im_a[5]_BAR ,
         \im_a[4]_BAR , \im_a[3]_BAR , \im_a[2]_BAR , \im_a[1]_BAR ,
         \im_a[0]_BAR ;
  wire   n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         \next_glb_cntr[1] , \next_write_addr_w[0] , \next_cr_y[0] , \h_1[2] ,
         \h_0[0] , \m_0[0] , \s_1[2] , \s_0[0] , N622, N623, N624, N625, N626,
         N627, N628, N629, N630, N631, N632, N633, N634, N635, N636, N637,
         N638, N639, N742, N743, N744, N745, N746, N747, N748, N750, N751,
         N752, N753, N754, N755, N756, N757, N758, N759, N760, N91, N92, N1453,
         N1454, N1455, N1456, N1457, N1458, N1459, N1460, N1667, N1668, N1669,
         N1670, N1671, N1672, N1673, N1674, N1675, N1676, N1677, N1678, N1679,
         N1680, N1681, N1682, N1683, N1684, N1685, N1686, N2282, N2283, N2284,
         N205, N2858, N2880, N2900, N2902, \C169/Z_0 , \C169/Z_1 , \C169/Z_2 ,
         \C169/Z_3 , \C169/Z_4 , \C169/Z_5 , \C169/Z_6 , \C169/Z_7 ,
         \C169/Z_8 , \C169/Z_9 , \C169/Z_10 , \C169/Z_11 , \C169/Z_12 ,
         \C169/Z_13 , \C169/Z_14 , \C169/Z_15 , \C169/Z_16 , \C169/Z_17 ,
         \C169/Z_18 , \C168/DATA3_0 , \C168/DATA3_1 , \C168/DATA3_2 ,
         \C168/DATA3_3 , \C168/DATA3_4 , \C168/DATA3_5 , \C168/DATA3_6 ,
         \C168/DATA3_7 , \C168/DATA3_8 , \C168/DATA3_9 , \C168/DATA3_10 ,
         \C168/DATA3_11 , \C168/DATA3_12 , \C168/DATA3_13 , \C168/DATA3_14 ,
         \C168/DATA3_15 , \C168/DATA3_16 , \C168/DATA3_17 , \C168/DATA3_18 ,
         \C168/DATA3_19 , n32, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n520, n521, n523, n524, n525, n526, n527, n528, n529,
         n530, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n545, n546, n547, n548, \DP_OP_719J1_125_1438/n26 ,
         \DP_OP_719J1_125_1438/n25 , \C1/Z_19 , \C1/Z_18 , \C1/Z_17 ,
         \C1/Z_16 , \C1/Z_15 , \C1/Z_14 , \C1/Z_13 , \C1/Z_12 , \C1/Z_11 ,
         \C1/Z_10 , \C1/Z_9 , \C1/Z_8 , \C1/Z_7 , \C1/Z_6 , \C1/Z_5 , \C1/Z_4 ,
         \U3/RSOP_717/C2/Z_19 , \U3/RSOP_717/C2/Z_18 , \U3/RSOP_717/C2/Z_17 ,
         \U3/RSOP_717/C2/Z_16 , \U3/RSOP_717/C2/Z_15 , \U3/RSOP_717/C2/Z_14 ,
         \U3/RSOP_717/C2/Z_13 , \U3/RSOP_717/C2/Z_12 , \U3/RSOP_717/C2/Z_11 ,
         \U3/RSOP_717/C2/Z_10 , \U3/RSOP_717/C2/Z_9 , \U3/RSOP_717/C2/Z_8 ,
         \U3/RSOP_717/C2/Z_7 , \U3/RSOP_717/C2/Z_6 , \U3/RSOP_717/C2/Z_5 ,
         \U3/RSOP_717/C2/Z_4 , \U3/RSOP_717/C2/Z_3 , \U3/RSOP_717/C2/Z_2 ,
         \U3/RSOP_717/C2/Z_1 , \U3/RSOP_717/C2/Z_0 , \C1/Z_3 , \C1/Z_2 ,
         \C1/Z_1 , \C1/Z_0 , \DP_OP_280J1_126_7605/I2 ,
         \DP_OP_280J1_126_7605/I3 , \DP_OP_280J1_126_7605/n27 ,
         \DP_OP_280J1_126_7605/n26 , \DP_OP_280J1_126_7605/n25 ,
         \DP_OP_280J1_126_7605/n24 , \DP_OP_280J1_126_7605/n23 ,
         \DP_OP_280J1_126_7605/n21 , \DP_OP_280J1_126_7605/n18 ,
         \DP_OP_280J1_126_7605/n17 , \DP_OP_280J1_126_7605/n16 ,
         \DP_OP_280J1_126_7605/n8 , \DP_OP_280J1_126_7605/n7 ,
         \DP_OP_280J1_126_7605/n6 , \DP_OP_280J1_126_7605/n5 ,
         \DP_OP_280J1_126_7605/n4 , \DP_OP_280J1_126_7605/n3 ,
         \DP_OP_280J1_126_7605/n2 , \DP_OP_280J1_126_7605/n1 ,
         \DP_OP_725J1_134_142/I2 , \DP_OP_725J1_134_142/I3 ,
         \DP_OP_725J1_134_142/I4 , \DP_OP_725J1_134_142/I7 ,
         \DP_OP_725J1_134_142/I10 , \DP_OP_725J1_134_142/n270 ,
         \DP_OP_725J1_134_142/n269 , \DP_OP_725J1_134_142/n268 ,
         \DP_OP_725J1_134_142/n267 , \DP_OP_725J1_134_142/n266 ,
         \DP_OP_725J1_134_142/n265 , \DP_OP_725J1_134_142/n264 ,
         \DP_OP_725J1_134_142/n263 , \DP_OP_725J1_134_142/n262 ,
         \DP_OP_725J1_134_142/n261 , \DP_OP_725J1_134_142/n260 ,
         \DP_OP_725J1_134_142/n259 , \DP_OP_725J1_134_142/n251 ,
         \DP_OP_725J1_134_142/n250 , \DP_OP_725J1_134_142/n249 ,
         \DP_OP_725J1_134_142/n248 , \DP_OP_725J1_134_142/n247 ,
         \DP_OP_725J1_134_142/n246 , \DP_OP_725J1_134_142/n245 ,
         \DP_OP_725J1_134_142/n244 , \DP_OP_725J1_134_142/n243 ,
         \DP_OP_725J1_134_142/n242 , \DP_OP_725J1_134_142/n241 ,
         \DP_OP_725J1_134_142/n240 , \DP_OP_725J1_134_142/n239 ,
         \DP_OP_725J1_134_142/n238 , \DP_OP_725J1_134_142/n237 ,
         \DP_OP_725J1_134_142/n236 , \DP_OP_725J1_134_142/n235 ,
         \DP_OP_725J1_134_142/n234 , \DP_OP_725J1_134_142/n233 ,
         \DP_OP_725J1_134_142/n232 , \DP_OP_725J1_134_142/n231 ,
         \DP_OP_725J1_134_142/n230 , \DP_OP_725J1_134_142/n229 ,
         \DP_OP_725J1_134_142/n228 , \DP_OP_725J1_134_142/n227 ,
         \DP_OP_725J1_134_142/n226 , \DP_OP_725J1_134_142/n225 ,
         \DP_OP_725J1_134_142/n224 , \DP_OP_725J1_134_142/n223 ,
         \DP_OP_725J1_134_142/n222 , \DP_OP_725J1_134_142/n221 ,
         \DP_OP_725J1_134_142/n220 , \DP_OP_725J1_134_142/n219 ,
         \DP_OP_725J1_134_142/n218 , \DP_OP_725J1_134_142/n217 ,
         \DP_OP_725J1_134_142/n216 , \DP_OP_725J1_134_142/n215 ,
         \DP_OP_725J1_134_142/n214 , \DP_OP_725J1_134_142/n213 ,
         \DP_OP_725J1_134_142/n206 , \DP_OP_725J1_134_142/n205 ,
         \DP_OP_725J1_134_142/n203 , \DP_OP_725J1_134_142/n202 ,
         \DP_OP_725J1_134_142/n200 , \DP_OP_725J1_134_142/n199 ,
         \DP_OP_725J1_134_142/n198 , \DP_OP_725J1_134_142/n197 ,
         \DP_OP_725J1_134_142/n196 , \DP_OP_725J1_134_142/n195 ,
         \DP_OP_725J1_134_142/n194 , \DP_OP_725J1_134_142/n193 ,
         \DP_OP_725J1_134_142/n192 , \DP_OP_725J1_134_142/n190 ,
         \DP_OP_725J1_134_142/n187 , \DP_OP_725J1_134_142/n184 ,
         \DP_OP_725J1_134_142/n183 , \DP_OP_725J1_134_142/n182 ,
         \DP_OP_725J1_134_142/n181 , \DP_OP_725J1_134_142/n180 ,
         \DP_OP_725J1_134_142/n179 , \DP_OP_725J1_134_142/n178 ,
         \DP_OP_725J1_134_142/n177 , \DP_OP_725J1_134_142/n176 ,
         \DP_OP_725J1_134_142/n175 , \DP_OP_725J1_134_142/n173 ,
         \DP_OP_725J1_134_142/n172 , \DP_OP_725J1_134_142/n171 ,
         \DP_OP_725J1_134_142/n170 , \DP_OP_725J1_134_142/n169 ,
         \DP_OP_725J1_134_142/n168 , \DP_OP_725J1_134_142/n167 ,
         \DP_OP_725J1_134_142/n166 , \DP_OP_725J1_134_142/n165 ,
         \DP_OP_725J1_134_142/n164 , \DP_OP_725J1_134_142/n163 ,
         \DP_OP_725J1_134_142/n162 , \DP_OP_725J1_134_142/n161 ,
         \DP_OP_725J1_134_142/n160 , \DP_OP_725J1_134_142/n159 ,
         \DP_OP_725J1_134_142/n158 , \DP_OP_725J1_134_142/n157 ,
         \DP_OP_725J1_134_142/n156 , \DP_OP_725J1_134_142/n155 ,
         \DP_OP_725J1_134_142/n154 , \DP_OP_725J1_134_142/n153 ,
         \DP_OP_725J1_134_142/n152 , \DP_OP_725J1_134_142/n151 ,
         \DP_OP_725J1_134_142/n150 , \DP_OP_725J1_134_142/n149 ,
         \DP_OP_725J1_134_142/n148 , \DP_OP_725J1_134_142/n147 ,
         \DP_OP_725J1_134_142/n146 , \DP_OP_725J1_134_142/n145 ,
         \DP_OP_725J1_134_142/n144 , \DP_OP_725J1_134_142/n143 ,
         \DP_OP_725J1_134_142/n142 , \DP_OP_725J1_134_142/n141 ,
         \DP_OP_725J1_134_142/n140 , \DP_OP_725J1_134_142/n138 ,
         \DP_OP_725J1_134_142/n137 , \DP_OP_725J1_134_142/n136 ,
         \DP_OP_725J1_134_142/n135 , \DP_OP_725J1_134_142/n134 ,
         \DP_OP_725J1_134_142/n133 , \DP_OP_725J1_134_142/n132 ,
         \DP_OP_725J1_134_142/n131 , \DP_OP_725J1_134_142/n130 ,
         \DP_OP_725J1_134_142/n129 , \DP_OP_725J1_134_142/n128 ,
         \DP_OP_725J1_134_142/n127 , \DP_OP_725J1_134_142/n126 ,
         \DP_OP_725J1_134_142/n125 , \DP_OP_725J1_134_142/n124 ,
         \DP_OP_725J1_134_142/n123 , \DP_OP_725J1_134_142/n122 ,
         \DP_OP_725J1_134_142/n121 , \DP_OP_725J1_134_142/n120 ,
         \DP_OP_725J1_134_142/n119 , \DP_OP_725J1_134_142/n118 ,
         \DP_OP_725J1_134_142/n117 , \DP_OP_725J1_134_142/n116 ,
         \DP_OP_725J1_134_142/n115 , \DP_OP_725J1_134_142/n114 ,
         \DP_OP_725J1_134_142/n113 , \DP_OP_725J1_134_142/n112 ,
         \DP_OP_725J1_134_142/n111 , \DP_OP_725J1_134_142/n110 ,
         \DP_OP_725J1_134_142/n109 , \DP_OP_725J1_134_142/n108 ,
         \DP_OP_725J1_134_142/n107 , \DP_OP_725J1_134_142/n106 ,
         \DP_OP_725J1_134_142/n105 , \DP_OP_725J1_134_142/n104 ,
         \DP_OP_725J1_134_142/n103 , \DP_OP_725J1_134_142/n102 ,
         \DP_OP_725J1_134_142/n101 , \DP_OP_725J1_134_142/n100 ,
         \DP_OP_725J1_134_142/n99 , \DP_OP_725J1_134_142/n98 ,
         \DP_OP_725J1_134_142/n97 , \DP_OP_725J1_134_142/n96 ,
         \DP_OP_725J1_134_142/n95 , \DP_OP_725J1_134_142/n94 ,
         \DP_OP_725J1_134_142/n93 , \DP_OP_725J1_134_142/n92 ,
         \DP_OP_725J1_134_142/n91 , \DP_OP_725J1_134_142/n90 ,
         \DP_OP_725J1_134_142/n89 , \DP_OP_725J1_134_142/n88 ,
         \DP_OP_725J1_134_142/n87 , \DP_OP_725J1_134_142/n86 ,
         \DP_OP_725J1_134_142/n85 , \DP_OP_725J1_134_142/n84 ,
         \DP_OP_725J1_134_142/n83 , \DP_OP_725J1_134_142/n82 ,
         \DP_OP_725J1_134_142/n81 , \DP_OP_725J1_134_142/n80 ,
         \DP_OP_725J1_134_142/n79 , \DP_OP_725J1_134_142/n78 ,
         \DP_OP_725J1_134_142/n77 , \DP_OP_725J1_134_142/n76 ,
         \DP_OP_725J1_134_142/n75 , \DP_OP_725J1_134_142/n74 ,
         \DP_OP_725J1_134_142/n73 , \DP_OP_725J1_134_142/n72 ,
         \DP_OP_725J1_134_142/n71 , \DP_OP_725J1_134_142/n70 ,
         \DP_OP_725J1_134_142/n69 , \DP_OP_725J1_134_142/n68 ,
         \DP_OP_725J1_134_142/n67 , \DP_OP_725J1_134_142/n66 ,
         \DP_OP_725J1_134_142/n65 , \DP_OP_725J1_134_142/n64 ,
         \DP_OP_725J1_134_142/n63 , \DP_OP_725J1_134_142/n62 ,
         \DP_OP_725J1_134_142/n61 , \DP_OP_725J1_134_142/n60 ,
         \DP_OP_725J1_134_142/n59 , \DP_OP_725J1_134_142/n58 ,
         \DP_OP_725J1_134_142/n57 , \DP_OP_725J1_134_142/n56 ,
         \DP_OP_725J1_134_142/n55 , \DP_OP_725J1_134_142/n54 ,
         \DP_OP_725J1_134_142/n53 , \DP_OP_725J1_134_142/n52 ,
         \DP_OP_725J1_134_142/n51 , \DP_OP_725J1_134_142/n50 ,
         \DP_OP_725J1_134_142/n49 , \DP_OP_725J1_134_142/n48 ,
         \DP_OP_725J1_134_142/n47 , \DP_OP_725J1_134_142/n46 ,
         \DP_OP_725J1_134_142/n45 , \DP_OP_725J1_134_142/n44 ,
         \DP_OP_725J1_134_142/n43 , \DP_OP_725J1_134_142/n42 ,
         \DP_OP_725J1_134_142/n41 , \DP_OP_725J1_134_142/n40 ,
         \DP_OP_725J1_134_142/n39 , \DP_OP_725J1_134_142/n38 ,
         \DP_OP_725J1_134_142/n37 , \DP_OP_725J1_134_142/n36 ,
         \DP_OP_725J1_134_142/n35 , \DP_OP_725J1_134_142/n34 ,
         \DP_OP_725J1_134_142/n33 , \DP_OP_725J1_134_142/n32 ,
         \DP_OP_725J1_134_142/n31 , \DP_OP_725J1_134_142/n30 ,
         \DP_OP_725J1_134_142/n29 , \DP_OP_725J1_134_142/n28 ,
         \DP_OP_725J1_134_142/n27 , \DP_OP_725J1_134_142/n26 ,
         \DP_OP_725J1_134_142/n25 , \DP_OP_725J1_134_142/n24 ,
         \DP_OP_725J1_134_142/n23 , \DP_OP_725J1_134_142/n22 ,
         \DP_OP_725J1_134_142/n21 , \DP_OP_725J1_134_142/n20 ,
         \DP_OP_725J1_134_142/n19 , \DP_OP_725J1_134_142/n18 ,
         \DP_OP_725J1_134_142/n17 , \DP_OP_725J1_134_142/n16 ,
         \DP_OP_725J1_134_142/n15 , \DP_OP_725J1_134_142/n14 ,
         \DP_OP_725J1_134_142/n13 , \DP_OP_725J1_134_142/n12 ,
         \DP_OP_725J1_134_142/n11 , \DP_OP_725J1_134_142/n10 ,
         \DP_OP_725J1_134_142/n9 , \DP_OP_725J1_134_142/n8 ,
         \DP_OP_725J1_134_142/n7 , \DP_OP_725J1_134_142/n6 ,
         \DP_OP_725J1_134_142/n5 , \DP_OP_725J1_134_142/n4 ,
         \DP_OP_725J1_134_142/n3 , \DP_OP_725J1_134_142/n2 ,
         \DP_OP_725J1_134_142/n1 , \intadd_3/A[8] , \intadd_3/A[7] ,
         \intadd_3/A[6] , \intadd_3/A[3] , \intadd_3/A[2] , \intadd_3/A[1] ,
         \intadd_3/A[0] , \intadd_3/B[6] , \intadd_3/B[5] , \intadd_3/B[4] ,
         \intadd_3/B[3] , \intadd_3/B[2] , \intadd_3/B[1] , \intadd_3/B[0] ,
         \intadd_3/CI , \intadd_3/SUM[8] , \intadd_3/SUM[7] ,
         \intadd_3/SUM[6] , \intadd_3/SUM[5] , \intadd_3/SUM[4] ,
         \intadd_3/SUM[3] , \intadd_3/SUM[2] , \intadd_3/SUM[1] ,
         \intadd_3/SUM[0] , \intadd_3/n9 , \intadd_3/n8 , \intadd_3/n7 ,
         \intadd_3/n6 , \intadd_3/n5 , \intadd_3/n4 , \intadd_3/n3 , n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n93, n95, n97, n99, n102, n103, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n211, n212,
         n213, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n522, n531, n532, n544, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971;
  wire   [2:0] next_state;
  wire   [2:0] state;
  wire   [19:0] work_cntr;
  wire   [19:0] next_work_cntr;
  wire   [19:0] global_cntr;
  wire   [19:0] write_addr;
  wire   [19:0] write_cntr;
  wire   [8:0] next_cr_x;
  wire   [3:0] m_1;
  wire   [19:0] read_cntr;
  wire   [8:0] cr_read_cntr;
  wire   [1:0] curr_photo;
  wire   [1:0] next_photo;
  assign \h_0[0]  = curr_time[16];
  assign \m_0[0]  = curr_time[8];
  assign \s_0[0]  = curr_time[0];
  assign en_init_time = N2858;
  assign en_curr_photo_addr = N2880;
  assign en_curr_photo_size = N2900;
  assign init_time_mux_sel = N2902;

  ADDHXL \DP_OP_280J1_126_7605/U16  ( .A(\C1/Z_0 ), .B(\C1/Z_1 ), .CO(
        \DP_OP_280J1_126_7605/n8 ), .S(\DP_OP_280J1_126_7605/n23 ) );
  ADDFXL \DP_OP_280J1_126_7605/U15  ( .A(\C1/Z_2 ), .B(\C1/Z_1 ), .CI(
        \DP_OP_280J1_126_7605/n8 ), .CO(\DP_OP_280J1_126_7605/n7 ), .S(
        \DP_OP_280J1_126_7605/n24 ) );
  ADDFXL \DP_OP_280J1_126_7605/U14  ( .A(\C1/Z_3 ), .B(\C1/Z_2 ), .CI(
        \DP_OP_280J1_126_7605/n7 ), .CO(\DP_OP_280J1_126_7605/n6 ), .S(
        \DP_OP_280J1_126_7605/n25 ) );
  ADDHXL \DP_OP_280J1_126_7605/U13  ( .A(\C1/Z_3 ), .B(
        \DP_OP_280J1_126_7605/n6 ), .CO(\DP_OP_280J1_126_7605/n27 ), .S(
        \DP_OP_280J1_126_7605/n26 ) );
  AO21X1 \DP_OP_280J1_126_7605/U11  ( .A0(\DP_OP_280J1_126_7605/n23 ), .A1(n85), .B0(\DP_OP_280J1_126_7605/I2 ), .Y(\DP_OP_280J1_126_7605/n17 ) );
  AO21X1 \DP_OP_280J1_126_7605/U10  ( .A0(\DP_OP_280J1_126_7605/n24 ), .A1(n85), .B0(\DP_OP_280J1_126_7605/I2 ), .Y(\DP_OP_280J1_126_7605/n18 ) );
  ADDHXL \DP_OP_725J1_134_142/U245  ( .A(write_addr[11]), .B(
        \DP_OP_725J1_134_142/n200 ), .CO(\DP_OP_725J1_134_142/n199 ), .S(
        \DP_OP_725J1_134_142/n261 ) );
  ADDHXL \DP_OP_725J1_134_142/U244  ( .A(n102), .B(\DP_OP_725J1_134_142/n199 ), 
        .CO(\DP_OP_725J1_134_142/n198 ), .S(\DP_OP_725J1_134_142/n262 ) );
  ADDHXL \DP_OP_725J1_134_142/U243  ( .A(n89), .B(\DP_OP_725J1_134_142/n198 ), 
        .CO(\DP_OP_725J1_134_142/n197 ), .S(\DP_OP_725J1_134_142/n263 ) );
  ADDHXL \DP_OP_725J1_134_142/U242  ( .A(n88), .B(\DP_OP_725J1_134_142/n197 ), 
        .CO(\DP_OP_725J1_134_142/n196 ), .S(\DP_OP_725J1_134_142/n264 ) );
  ADDHXL \DP_OP_725J1_134_142/U241  ( .A(write_addr[15]), .B(
        \DP_OP_725J1_134_142/n196 ), .CO(\DP_OP_725J1_134_142/n195 ), .S(
        \DP_OP_725J1_134_142/n265 ) );
  ADDHXL \DP_OP_725J1_134_142/U240  ( .A(write_addr[16]), .B(
        \DP_OP_725J1_134_142/n195 ), .CO(\DP_OP_725J1_134_142/n194 ), .S(
        \DP_OP_725J1_134_142/n266 ) );
  ADDHXL \DP_OP_725J1_134_142/U239  ( .A(write_addr[17]), .B(
        \DP_OP_725J1_134_142/n194 ), .CO(\DP_OP_725J1_134_142/n193 ), .S(
        \DP_OP_725J1_134_142/n267 ) );
  ADDHXL \DP_OP_725J1_134_142/U238  ( .A(write_addr[18]), .B(
        \DP_OP_725J1_134_142/n193 ), .CO(\DP_OP_725J1_134_142/n192 ), .S(
        \DP_OP_725J1_134_142/n268 ) );
  ADDHXL \DP_OP_725J1_134_142/U237  ( .A(write_addr[19]), .B(
        \DP_OP_725J1_134_142/n192 ), .CO(\DP_OP_725J1_134_142/n270 ), .S(
        \DP_OP_725J1_134_142/n269 ) );
  ADDHXL \DP_OP_725J1_134_142/U223  ( .A(n88), .B(\DP_OP_725J1_134_142/n180 ), 
        .CO(\DP_OP_725J1_134_142/n179 ), .S(N633) );
  ADDFXL \DP_OP_725J1_134_142/U204  ( .A(N742), .B(fb_addr[1]), .CI(
        \DP_OP_725J1_134_142/n164 ), .CO(\DP_OP_725J1_134_142/n163 ), .S(N1668) );
  ADDFXL \DP_OP_725J1_134_142/U203  ( .A(N743), .B(fb_addr[2]), .CI(
        \DP_OP_725J1_134_142/n163 ), .CO(\DP_OP_725J1_134_142/n162 ), .S(N1669) );
  ADDFXL \DP_OP_725J1_134_142/U202  ( .A(N744), .B(fb_addr[3]), .CI(
        \DP_OP_725J1_134_142/n162 ), .CO(\DP_OP_725J1_134_142/n161 ), .S(N1670) );
  ADDFXL \DP_OP_725J1_134_142/U201  ( .A(N745), .B(fb_addr[4]), .CI(
        \DP_OP_725J1_134_142/n161 ), .CO(\DP_OP_725J1_134_142/n160 ), .S(N1671) );
  ADDFXL \DP_OP_725J1_134_142/U200  ( .A(N746), .B(fb_addr[5]), .CI(
        \DP_OP_725J1_134_142/n160 ), .CO(\DP_OP_725J1_134_142/n159 ), .S(N1672) );
  ADDFXL \DP_OP_725J1_134_142/U199  ( .A(N747), .B(fb_addr[6]), .CI(
        \DP_OP_725J1_134_142/n159 ), .CO(\DP_OP_725J1_134_142/n158 ), .S(N1673) );
  ADDFXL \DP_OP_725J1_134_142/U198  ( .A(N748), .B(fb_addr[7]), .CI(
        \DP_OP_725J1_134_142/n158 ), .CO(\DP_OP_725J1_134_142/n157 ), .S(N1674) );
  ADDFXL \DP_OP_725J1_134_142/U197  ( .A(write_addr[8]), .B(fb_addr[8]), .CI(
        \DP_OP_725J1_134_142/n157 ), .CO(\DP_OP_725J1_134_142/n156 ), .S(N1675) );
  ADDFXL \DP_OP_725J1_134_142/U196  ( .A(write_addr[9]), .B(fb_addr[9]), .CI(
        \DP_OP_725J1_134_142/n156 ), .CO(\DP_OP_725J1_134_142/n155 ), .S(N1676) );
  ADDFXL \DP_OP_725J1_134_142/U195  ( .A(write_addr[10]), .B(fb_addr[10]), 
        .CI(\DP_OP_725J1_134_142/n155 ), .CO(\DP_OP_725J1_134_142/n154 ), .S(
        N1677) );
  ADDFXL \DP_OP_725J1_134_142/U194  ( .A(write_addr[11]), .B(fb_addr[11]), 
        .CI(\DP_OP_725J1_134_142/n154 ), .CO(\DP_OP_725J1_134_142/n153 ), .S(
        N1678) );
  ADDFXL \DP_OP_725J1_134_142/U193  ( .A(n102), .B(fb_addr[12]), .CI(
        \DP_OP_725J1_134_142/n153 ), .CO(\DP_OP_725J1_134_142/n152 ), .S(N1679) );
  ADDFXL \DP_OP_725J1_134_142/U192  ( .A(n89), .B(fb_addr[13]), .CI(
        \DP_OP_725J1_134_142/n152 ), .CO(\DP_OP_725J1_134_142/n151 ), .S(N1680) );
  ADDFXL \DP_OP_725J1_134_142/U191  ( .A(n88), .B(fb_addr[14]), .CI(
        \DP_OP_725J1_134_142/n151 ), .CO(\DP_OP_725J1_134_142/n150 ), .S(N1681) );
  ADDFXL \DP_OP_725J1_134_142/U190  ( .A(write_addr[15]), .B(fb_addr[15]), 
        .CI(\DP_OP_725J1_134_142/n150 ), .CO(\DP_OP_725J1_134_142/n149 ), .S(
        N1682) );
  ADDFXL \DP_OP_725J1_134_142/U189  ( .A(write_addr[16]), .B(fb_addr[16]), 
        .CI(\DP_OP_725J1_134_142/n149 ), .CO(\DP_OP_725J1_134_142/n148 ), .S(
        N1683) );
  ADDFXL \DP_OP_725J1_134_142/U188  ( .A(write_addr[17]), .B(fb_addr[17]), 
        .CI(\DP_OP_725J1_134_142/n148 ), .CO(\DP_OP_725J1_134_142/n147 ), .S(
        N1684) );
  ADDFXL \DP_OP_725J1_134_142/U187  ( .A(write_addr[18]), .B(fb_addr[18]), 
        .CI(\DP_OP_725J1_134_142/n147 ), .CO(\DP_OP_725J1_134_142/n146 ), .S(
        N1685) );
  AO22X1 \DP_OP_725J1_134_142/U22  ( .A0(N1686), .A1(si_sel), .B0(
        \DP_OP_725J1_134_142/I10 ), .B1(\U3/RSOP_717/C2/Z_19 ), .Y(
        \DP_OP_725J1_134_142/n232 ) );
  ADDHXL \DP_OP_725J1_134_142/U21  ( .A(n761), .B(\DP_OP_725J1_134_142/n213 ), 
        .CO(\DP_OP_725J1_134_142/n20 ), .S(\C168/DATA3_0 ) );
  ADDFXL \DP_OP_725J1_134_142/U20  ( .A(\DP_OP_725J1_134_142/n20 ), .B(n762), 
        .CI(\DP_OP_725J1_134_142/n214 ), .CO(\DP_OP_725J1_134_142/n19 ), .S(
        \C168/DATA3_1 ) );
  ADDFXL \DP_OP_725J1_134_142/U19  ( .A(\DP_OP_725J1_134_142/n215 ), .B(n763), 
        .CI(\DP_OP_725J1_134_142/n19 ), .CO(\DP_OP_725J1_134_142/n18 ), .S(
        \C168/DATA3_2 ) );
  ADDFXL \DP_OP_725J1_134_142/U18  ( .A(\DP_OP_725J1_134_142/n216 ), .B(n764), 
        .CI(\DP_OP_725J1_134_142/n18 ), .CO(\DP_OP_725J1_134_142/n17 ), .S(
        \C168/DATA3_3 ) );
  ADDFXL \DP_OP_725J1_134_142/U17  ( .A(\DP_OP_725J1_134_142/n217 ), .B(
        \C1/Z_4 ), .CI(\DP_OP_725J1_134_142/n17 ), .CO(
        \DP_OP_725J1_134_142/n16 ), .S(\C168/DATA3_4 ) );
  ADDFXL \DP_OP_725J1_134_142/U16  ( .A(\DP_OP_725J1_134_142/n218 ), .B(
        \C1/Z_5 ), .CI(\DP_OP_725J1_134_142/n16 ), .CO(
        \DP_OP_725J1_134_142/n15 ), .S(\C168/DATA3_5 ) );
  ADDFXL \DP_OP_725J1_134_142/U15  ( .A(\DP_OP_725J1_134_142/n219 ), .B(
        \C1/Z_6 ), .CI(\DP_OP_725J1_134_142/n15 ), .CO(
        \DP_OP_725J1_134_142/n14 ), .S(\C168/DATA3_6 ) );
  ADDFXL \DP_OP_725J1_134_142/U14  ( .A(\DP_OP_725J1_134_142/n220 ), .B(
        \C1/Z_7 ), .CI(\DP_OP_725J1_134_142/n14 ), .CO(
        \DP_OP_725J1_134_142/n13 ), .S(\C168/DATA3_7 ) );
  ADDFXL \DP_OP_725J1_134_142/U13  ( .A(\DP_OP_725J1_134_142/n221 ), .B(
        \C1/Z_8 ), .CI(\DP_OP_725J1_134_142/n13 ), .CO(
        \DP_OP_725J1_134_142/n12 ), .S(\C168/DATA3_8 ) );
  ADDFXL \DP_OP_725J1_134_142/U12  ( .A(\DP_OP_725J1_134_142/n222 ), .B(
        \C1/Z_9 ), .CI(\DP_OP_725J1_134_142/n12 ), .CO(
        \DP_OP_725J1_134_142/n11 ), .S(\C168/DATA3_9 ) );
  ADDFXL \DP_OP_725J1_134_142/U11  ( .A(\DP_OP_725J1_134_142/n223 ), .B(
        \C1/Z_10 ), .CI(\DP_OP_725J1_134_142/n11 ), .CO(
        \DP_OP_725J1_134_142/n10 ), .S(\C168/DATA3_10 ) );
  ADDFXL \DP_OP_725J1_134_142/U10  ( .A(\DP_OP_725J1_134_142/n224 ), .B(
        \C1/Z_11 ), .CI(\DP_OP_725J1_134_142/n10 ), .CO(
        \DP_OP_725J1_134_142/n9 ), .S(\C168/DATA3_11 ) );
  ADDFXL \DP_OP_725J1_134_142/U9  ( .A(\DP_OP_725J1_134_142/n225 ), .B(
        \C1/Z_12 ), .CI(\DP_OP_725J1_134_142/n9 ), .CO(
        \DP_OP_725J1_134_142/n8 ), .S(\C168/DATA3_12 ) );
  ADDFXL \DP_OP_725J1_134_142/U8  ( .A(\DP_OP_725J1_134_142/n226 ), .B(
        \C1/Z_13 ), .CI(\DP_OP_725J1_134_142/n8 ), .CO(
        \DP_OP_725J1_134_142/n7 ), .S(\C168/DATA3_13 ) );
  ADDFXL \DP_OP_725J1_134_142/U7  ( .A(\DP_OP_725J1_134_142/n227 ), .B(
        \C1/Z_14 ), .CI(\DP_OP_725J1_134_142/n7 ), .CO(
        \DP_OP_725J1_134_142/n6 ), .S(\C168/DATA3_14 ) );
  ADDFXL \DP_OP_725J1_134_142/U6  ( .A(\DP_OP_725J1_134_142/n228 ), .B(
        \C1/Z_15 ), .CI(\DP_OP_725J1_134_142/n6 ), .CO(
        \DP_OP_725J1_134_142/n5 ), .S(\C168/DATA3_15 ) );
  ADDFXL \DP_OP_725J1_134_142/U5  ( .A(\DP_OP_725J1_134_142/n229 ), .B(
        \C1/Z_16 ), .CI(\DP_OP_725J1_134_142/n5 ), .CO(
        \DP_OP_725J1_134_142/n4 ), .S(\C168/DATA3_16 ) );
  ADDFXL \DP_OP_725J1_134_142/U4  ( .A(\DP_OP_725J1_134_142/n230 ), .B(
        \C1/Z_17 ), .CI(\DP_OP_725J1_134_142/n4 ), .CO(
        \DP_OP_725J1_134_142/n3 ), .S(\C168/DATA3_17 ) );
  ADDFXL \DP_OP_725J1_134_142/U3  ( .A(\DP_OP_725J1_134_142/n231 ), .B(
        \C1/Z_18 ), .CI(\DP_OP_725J1_134_142/n3 ), .CO(
        \DP_OP_725J1_134_142/n2 ), .S(\C168/DATA3_18 ) );
  ADDFXL \intadd_3/U10  ( .A(\intadd_3/A[0] ), .B(\intadd_3/B[0] ), .CI(
        \intadd_3/CI ), .CO(\intadd_3/n9 ), .S(\intadd_3/SUM[0] ) );
  ADDFXL \intadd_3/U9  ( .A(\intadd_3/A[1] ), .B(\intadd_3/B[1] ), .CI(
        \intadd_3/n9 ), .CO(\intadd_3/n8 ), .S(\intadd_3/SUM[1] ) );
  ADDFXL \intadd_3/U8  ( .A(\intadd_3/A[2] ), .B(\intadd_3/B[2] ), .CI(
        \intadd_3/n8 ), .CO(\intadd_3/n7 ), .S(\intadd_3/SUM[2] ) );
  ADDFXL \intadd_3/U7  ( .A(\intadd_3/A[3] ), .B(\intadd_3/B[3] ), .CI(
        \intadd_3/n7 ), .CO(\intadd_3/n6 ), .S(\intadd_3/SUM[3] ) );
  ADDFXL \intadd_3/U6  ( .A(\DP_OP_719J1_125_1438/n26 ), .B(\intadd_3/B[4] ), 
        .CI(\intadd_3/n6 ), .CO(\intadd_3/n5 ), .S(\intadd_3/SUM[4] ) );
  ADDFXL \intadd_3/U5  ( .A(\DP_OP_719J1_125_1438/n25 ), .B(\intadd_3/B[5] ), 
        .CI(\intadd_3/n5 ), .CO(\intadd_3/n4 ), .S(\intadd_3/SUM[5] ) );
  ADDFXL \intadd_3/U4  ( .A(\intadd_3/A[6] ), .B(\intadd_3/B[6] ), .CI(
        \intadd_3/n4 ), .CO(\intadd_3/n3 ), .S(\intadd_3/SUM[6] ) );
  DFFRX1 \cr_read_cntr_reg/q_reg[7]  ( .D(n495), .CK(clk), .RN(n43), .QN(n237)
         );
  DFFRX1 \cr_read_cntr_reg/q_reg[8]  ( .D(n494), .CK(clk), .RN(n43), .Q(
        cr_read_cntr[8]) );
  NAND2X1 \DP_OP_725J1_134_142/U101  ( .A(N639), .B(\DP_OP_725J1_134_142/I2 ), 
        .Y(\DP_OP_725J1_134_142/n79 ) );
  NAND2X1 \DP_OP_725J1_134_142/U106  ( .A(N638), .B(\DP_OP_725J1_134_142/I2 ), 
        .Y(\DP_OP_725J1_134_142/n83 ) );
  NAND2X1 \DP_OP_725J1_134_142/U111  ( .A(N637), .B(\DP_OP_725J1_134_142/I2 ), 
        .Y(\DP_OP_725J1_134_142/n87 ) );
  NAND2X1 \DP_OP_725J1_134_142/U116  ( .A(N636), .B(\DP_OP_725J1_134_142/I2 ), 
        .Y(\DP_OP_725J1_134_142/n91 ) );
  NAND2X1 \DP_OP_725J1_134_142/U121  ( .A(N635), .B(\DP_OP_725J1_134_142/I2 ), 
        .Y(\DP_OP_725J1_134_142/n95 ) );
  NAND2X1 \DP_OP_725J1_134_142/U126  ( .A(N634), .B(\DP_OP_725J1_134_142/I2 ), 
        .Y(\DP_OP_725J1_134_142/n99 ) );
  NAND2X1 \DP_OP_725J1_134_142/U131  ( .A(n57), .B(\DP_OP_725J1_134_142/I2 ), 
        .Y(\DP_OP_725J1_134_142/n103 ) );
  NAND2X1 \DP_OP_725J1_134_142/U136  ( .A(N632), .B(\DP_OP_725J1_134_142/I2 ), 
        .Y(\DP_OP_725J1_134_142/n107 ) );
  NAND2X1 \DP_OP_725J1_134_142/U141  ( .A(N631), .B(\DP_OP_725J1_134_142/I2 ), 
        .Y(\DP_OP_725J1_134_142/n111 ) );
  NAND2X1 \DP_OP_725J1_134_142/U146  ( .A(N630), .B(\DP_OP_725J1_134_142/I2 ), 
        .Y(\DP_OP_725J1_134_142/n115 ) );
  NAND2X1 \DP_OP_725J1_134_142/U151  ( .A(N629), .B(\DP_OP_725J1_134_142/I2 ), 
        .Y(\DP_OP_725J1_134_142/n119 ) );
  NAND2X1 \DP_OP_725J1_134_142/U155  ( .A(N628), .B(\DP_OP_725J1_134_142/I2 ), 
        .Y(\DP_OP_725J1_134_142/n122 ) );
  AOI22X1 \DP_OP_725J1_134_142/U157  ( .A0(n233), .A1(\DP_OP_725J1_134_142/I4 ), .B0(n209), .B1(\C169/Z_7 ), .Y(\DP_OP_725J1_134_142/n124 ) );
  NAND2X1 \DP_OP_725J1_134_142/U160  ( .A(N627), .B(\DP_OP_725J1_134_142/I2 ), 
        .Y(\DP_OP_725J1_134_142/n126 ) );
  AOI22X1 \DP_OP_725J1_134_142/U161  ( .A0(n209), .A1(\C169/Z_6 ), .B0(
        \DP_OP_725J1_134_142/I4 ), .B1(N748), .Y(\DP_OP_725J1_134_142/n127 )
         );
  ADDHXL \DP_OP_280J1_126_7605/U6  ( .A(N91), .B(\DP_OP_280J1_126_7605/n16 ), 
        .CO(\DP_OP_280J1_126_7605/n5 ), .S(N1456) );
  ADDFXL \DP_OP_280J1_126_7605/U5  ( .A(\DP_OP_280J1_126_7605/n5 ), .B(N92), 
        .CI(\DP_OP_280J1_126_7605/n17 ), .CO(\DP_OP_280J1_126_7605/n4 ), .S(
        N1457) );
  ADDHXL \DP_OP_280J1_126_7605/U4  ( .A(\DP_OP_280J1_126_7605/n4 ), .B(
        \DP_OP_280J1_126_7605/n18 ), .CO(\DP_OP_280J1_126_7605/n3 ), .S(N1458)
         );
  NAND2XL \DP_OP_725J1_134_142/U24  ( .A(N1685), .B(si_sel), .Y(
        \DP_OP_725J1_134_142/n21 ) );
  NAND2XL \DP_OP_725J1_134_142/U100  ( .A(\DP_OP_725J1_134_142/n270 ), .B(
        \DP_OP_725J1_134_142/I3 ), .Y(\DP_OP_725J1_134_142/n78 ) );
  NAND2XL \DP_OP_725J1_134_142/U102  ( .A(N760), .B(\DP_OP_725J1_134_142/I4 ), 
        .Y(\DP_OP_725J1_134_142/n80 ) );
  NAND2XL \DP_OP_725J1_134_142/U103  ( .A(n209), .B(\C169/Z_18 ), .Y(
        \DP_OP_725J1_134_142/n81 ) );
  NAND4XL \DP_OP_725J1_134_142/U99  ( .A(\DP_OP_725J1_134_142/n78 ), .B(
        \DP_OP_725J1_134_142/n79 ), .C(\DP_OP_725J1_134_142/n80 ), .D(
        \DP_OP_725J1_134_142/n81 ), .Y(\DP_OP_725J1_134_142/n251 ) );
  NAND2XL \DP_OP_725J1_134_142/U25  ( .A(\DP_OP_725J1_134_142/n251 ), .B(
        \DP_OP_725J1_134_142/I7 ), .Y(\DP_OP_725J1_134_142/n22 ) );
  NAND2XL \DP_OP_725J1_134_142/U26  ( .A(\DP_OP_725J1_134_142/I10 ), .B(
        \U3/RSOP_717/C2/Z_18 ), .Y(\DP_OP_725J1_134_142/n23 ) );
  NAND3XL \DP_OP_725J1_134_142/U23  ( .A(\DP_OP_725J1_134_142/n21 ), .B(
        \DP_OP_725J1_134_142/n22 ), .C(\DP_OP_725J1_134_142/n23 ), .Y(
        \DP_OP_725J1_134_142/n231 ) );
  NAND2XL \DP_OP_725J1_134_142/U28  ( .A(N1684), .B(si_sel), .Y(
        \DP_OP_725J1_134_142/n24 ) );
  NAND2XL \DP_OP_725J1_134_142/U105  ( .A(\DP_OP_725J1_134_142/n269 ), .B(
        \DP_OP_725J1_134_142/I3 ), .Y(\DP_OP_725J1_134_142/n82 ) );
  NAND2XL \DP_OP_725J1_134_142/U107  ( .A(N759), .B(\DP_OP_725J1_134_142/I4 ), 
        .Y(\DP_OP_725J1_134_142/n84 ) );
  NAND2XL \DP_OP_725J1_134_142/U108  ( .A(n209), .B(\C169/Z_17 ), .Y(
        \DP_OP_725J1_134_142/n85 ) );
  NAND4XL \DP_OP_725J1_134_142/U104  ( .A(\DP_OP_725J1_134_142/n82 ), .B(
        \DP_OP_725J1_134_142/n83 ), .C(\DP_OP_725J1_134_142/n84 ), .D(
        \DP_OP_725J1_134_142/n85 ), .Y(\DP_OP_725J1_134_142/n250 ) );
  NAND2XL \DP_OP_725J1_134_142/U29  ( .A(\DP_OP_725J1_134_142/n250 ), .B(
        \DP_OP_725J1_134_142/I7 ), .Y(\DP_OP_725J1_134_142/n25 ) );
  NAND2XL \DP_OP_725J1_134_142/U30  ( .A(\DP_OP_725J1_134_142/I10 ), .B(
        \U3/RSOP_717/C2/Z_17 ), .Y(\DP_OP_725J1_134_142/n26 ) );
  NAND3XL \DP_OP_725J1_134_142/U27  ( .A(\DP_OP_725J1_134_142/n24 ), .B(
        \DP_OP_725J1_134_142/n25 ), .C(\DP_OP_725J1_134_142/n26 ), .Y(
        \DP_OP_725J1_134_142/n230 ) );
  NAND2XL \DP_OP_725J1_134_142/U32  ( .A(N1683), .B(si_sel), .Y(
        \DP_OP_725J1_134_142/n27 ) );
  NAND2XL \DP_OP_725J1_134_142/U110  ( .A(\DP_OP_725J1_134_142/n268 ), .B(
        \DP_OP_725J1_134_142/I3 ), .Y(\DP_OP_725J1_134_142/n86 ) );
  NAND2XL \DP_OP_725J1_134_142/U112  ( .A(N758), .B(\DP_OP_725J1_134_142/I4 ), 
        .Y(\DP_OP_725J1_134_142/n88 ) );
  NAND2XL \DP_OP_725J1_134_142/U113  ( .A(n209), .B(\C169/Z_16 ), .Y(
        \DP_OP_725J1_134_142/n89 ) );
  NAND4XL \DP_OP_725J1_134_142/U109  ( .A(\DP_OP_725J1_134_142/n86 ), .B(
        \DP_OP_725J1_134_142/n87 ), .C(\DP_OP_725J1_134_142/n88 ), .D(
        \DP_OP_725J1_134_142/n89 ), .Y(\DP_OP_725J1_134_142/n249 ) );
  NAND2XL \DP_OP_725J1_134_142/U33  ( .A(\DP_OP_725J1_134_142/n249 ), .B(
        \DP_OP_725J1_134_142/I7 ), .Y(\DP_OP_725J1_134_142/n28 ) );
  NAND2XL \DP_OP_725J1_134_142/U34  ( .A(\DP_OP_725J1_134_142/I10 ), .B(
        \U3/RSOP_717/C2/Z_16 ), .Y(\DP_OP_725J1_134_142/n29 ) );
  NAND3XL \DP_OP_725J1_134_142/U31  ( .A(\DP_OP_725J1_134_142/n27 ), .B(
        \DP_OP_725J1_134_142/n28 ), .C(\DP_OP_725J1_134_142/n29 ), .Y(
        \DP_OP_725J1_134_142/n229 ) );
  NAND2XL \DP_OP_725J1_134_142/U36  ( .A(N1682), .B(si_sel), .Y(
        \DP_OP_725J1_134_142/n30 ) );
  NAND2XL \DP_OP_725J1_134_142/U115  ( .A(\DP_OP_725J1_134_142/n267 ), .B(
        \DP_OP_725J1_134_142/I3 ), .Y(\DP_OP_725J1_134_142/n90 ) );
  NAND2XL \DP_OP_725J1_134_142/U117  ( .A(N757), .B(\DP_OP_725J1_134_142/I4 ), 
        .Y(\DP_OP_725J1_134_142/n92 ) );
  NAND2XL \DP_OP_725J1_134_142/U118  ( .A(n209), .B(\C169/Z_15 ), .Y(
        \DP_OP_725J1_134_142/n93 ) );
  NAND4XL \DP_OP_725J1_134_142/U114  ( .A(\DP_OP_725J1_134_142/n90 ), .B(
        \DP_OP_725J1_134_142/n91 ), .C(\DP_OP_725J1_134_142/n92 ), .D(
        \DP_OP_725J1_134_142/n93 ), .Y(\DP_OP_725J1_134_142/n248 ) );
  NAND2XL \DP_OP_725J1_134_142/U37  ( .A(\DP_OP_725J1_134_142/n248 ), .B(
        \DP_OP_725J1_134_142/I7 ), .Y(\DP_OP_725J1_134_142/n31 ) );
  NAND2XL \DP_OP_725J1_134_142/U38  ( .A(\DP_OP_725J1_134_142/I10 ), .B(
        \U3/RSOP_717/C2/Z_15 ), .Y(\DP_OP_725J1_134_142/n32 ) );
  NAND3XL \DP_OP_725J1_134_142/U35  ( .A(\DP_OP_725J1_134_142/n30 ), .B(
        \DP_OP_725J1_134_142/n31 ), .C(\DP_OP_725J1_134_142/n32 ), .Y(
        \DP_OP_725J1_134_142/n228 ) );
  NAND2XL \DP_OP_725J1_134_142/U40  ( .A(N1681), .B(si_sel), .Y(
        \DP_OP_725J1_134_142/n33 ) );
  NAND2XL \DP_OP_725J1_134_142/U120  ( .A(\DP_OP_725J1_134_142/n266 ), .B(
        \DP_OP_725J1_134_142/I3 ), .Y(\DP_OP_725J1_134_142/n94 ) );
  NAND2XL \DP_OP_725J1_134_142/U122  ( .A(N756), .B(\DP_OP_725J1_134_142/I4 ), 
        .Y(\DP_OP_725J1_134_142/n96 ) );
  NAND2XL \DP_OP_725J1_134_142/U123  ( .A(n209), .B(\C169/Z_14 ), .Y(
        \DP_OP_725J1_134_142/n97 ) );
  NAND4XL \DP_OP_725J1_134_142/U119  ( .A(\DP_OP_725J1_134_142/n94 ), .B(
        \DP_OP_725J1_134_142/n95 ), .C(\DP_OP_725J1_134_142/n96 ), .D(
        \DP_OP_725J1_134_142/n97 ), .Y(\DP_OP_725J1_134_142/n247 ) );
  NAND2XL \DP_OP_725J1_134_142/U41  ( .A(\DP_OP_725J1_134_142/n247 ), .B(
        \DP_OP_725J1_134_142/I7 ), .Y(\DP_OP_725J1_134_142/n34 ) );
  NAND2XL \DP_OP_725J1_134_142/U42  ( .A(\DP_OP_725J1_134_142/I10 ), .B(
        \U3/RSOP_717/C2/Z_14 ), .Y(\DP_OP_725J1_134_142/n35 ) );
  NAND3XL \DP_OP_725J1_134_142/U39  ( .A(\DP_OP_725J1_134_142/n33 ), .B(
        \DP_OP_725J1_134_142/n34 ), .C(\DP_OP_725J1_134_142/n35 ), .Y(
        \DP_OP_725J1_134_142/n227 ) );
  NAND2XL \DP_OP_725J1_134_142/U44  ( .A(N1680), .B(si_sel), .Y(
        \DP_OP_725J1_134_142/n36 ) );
  NAND2XL \DP_OP_725J1_134_142/U125  ( .A(\DP_OP_725J1_134_142/n265 ), .B(
        \DP_OP_725J1_134_142/I3 ), .Y(\DP_OP_725J1_134_142/n98 ) );
  NAND2XL \DP_OP_725J1_134_142/U127  ( .A(N755), .B(\DP_OP_725J1_134_142/I4 ), 
        .Y(\DP_OP_725J1_134_142/n100 ) );
  NAND2XL \DP_OP_725J1_134_142/U128  ( .A(n209), .B(\C169/Z_13 ), .Y(
        \DP_OP_725J1_134_142/n101 ) );
  NAND4XL \DP_OP_725J1_134_142/U124  ( .A(\DP_OP_725J1_134_142/n98 ), .B(
        \DP_OP_725J1_134_142/n99 ), .C(\DP_OP_725J1_134_142/n100 ), .D(
        \DP_OP_725J1_134_142/n101 ), .Y(\DP_OP_725J1_134_142/n246 ) );
  NAND2XL \DP_OP_725J1_134_142/U45  ( .A(\DP_OP_725J1_134_142/n246 ), .B(
        \DP_OP_725J1_134_142/I7 ), .Y(\DP_OP_725J1_134_142/n37 ) );
  NAND2XL \DP_OP_725J1_134_142/U46  ( .A(\DP_OP_725J1_134_142/I10 ), .B(
        \U3/RSOP_717/C2/Z_13 ), .Y(\DP_OP_725J1_134_142/n38 ) );
  NAND3XL \DP_OP_725J1_134_142/U43  ( .A(\DP_OP_725J1_134_142/n36 ), .B(
        \DP_OP_725J1_134_142/n37 ), .C(\DP_OP_725J1_134_142/n38 ), .Y(
        \DP_OP_725J1_134_142/n226 ) );
  NAND2XL \DP_OP_725J1_134_142/U48  ( .A(N1679), .B(si_sel), .Y(
        \DP_OP_725J1_134_142/n39 ) );
  NAND2XL \DP_OP_725J1_134_142/U130  ( .A(\DP_OP_725J1_134_142/n264 ), .B(
        \DP_OP_725J1_134_142/I3 ), .Y(\DP_OP_725J1_134_142/n102 ) );
  NAND2XL \DP_OP_725J1_134_142/U132  ( .A(N754), .B(\DP_OP_725J1_134_142/I4 ), 
        .Y(\DP_OP_725J1_134_142/n104 ) );
  NAND2XL \DP_OP_725J1_134_142/U133  ( .A(n209), .B(\C169/Z_12 ), .Y(
        \DP_OP_725J1_134_142/n105 ) );
  NAND4XL \DP_OP_725J1_134_142/U129  ( .A(\DP_OP_725J1_134_142/n102 ), .B(
        \DP_OP_725J1_134_142/n103 ), .C(\DP_OP_725J1_134_142/n104 ), .D(
        \DP_OP_725J1_134_142/n105 ), .Y(\DP_OP_725J1_134_142/n245 ) );
  NAND2XL \DP_OP_725J1_134_142/U49  ( .A(\DP_OP_725J1_134_142/n245 ), .B(
        \DP_OP_725J1_134_142/I7 ), .Y(\DP_OP_725J1_134_142/n40 ) );
  NAND2XL \DP_OP_725J1_134_142/U50  ( .A(\DP_OP_725J1_134_142/I10 ), .B(
        \U3/RSOP_717/C2/Z_12 ), .Y(\DP_OP_725J1_134_142/n41 ) );
  NAND3XL \DP_OP_725J1_134_142/U47  ( .A(\DP_OP_725J1_134_142/n39 ), .B(
        \DP_OP_725J1_134_142/n40 ), .C(\DP_OP_725J1_134_142/n41 ), .Y(
        \DP_OP_725J1_134_142/n225 ) );
  NAND2XL \DP_OP_725J1_134_142/U52  ( .A(N1678), .B(si_sel), .Y(
        \DP_OP_725J1_134_142/n42 ) );
  NAND2XL \DP_OP_725J1_134_142/U135  ( .A(\DP_OP_725J1_134_142/n263 ), .B(
        \DP_OP_725J1_134_142/I3 ), .Y(\DP_OP_725J1_134_142/n106 ) );
  NAND2XL \DP_OP_725J1_134_142/U137  ( .A(N753), .B(\DP_OP_725J1_134_142/I4 ), 
        .Y(\DP_OP_725J1_134_142/n108 ) );
  NAND2XL \DP_OP_725J1_134_142/U138  ( .A(n209), .B(\C169/Z_11 ), .Y(
        \DP_OP_725J1_134_142/n109 ) );
  NAND4XL \DP_OP_725J1_134_142/U134  ( .A(\DP_OP_725J1_134_142/n106 ), .B(
        \DP_OP_725J1_134_142/n107 ), .C(\DP_OP_725J1_134_142/n108 ), .D(
        \DP_OP_725J1_134_142/n109 ), .Y(\DP_OP_725J1_134_142/n244 ) );
  NAND2XL \DP_OP_725J1_134_142/U53  ( .A(\DP_OP_725J1_134_142/n244 ), .B(
        \DP_OP_725J1_134_142/I7 ), .Y(\DP_OP_725J1_134_142/n43 ) );
  NAND2XL \DP_OP_725J1_134_142/U54  ( .A(\DP_OP_725J1_134_142/I10 ), .B(
        \U3/RSOP_717/C2/Z_11 ), .Y(\DP_OP_725J1_134_142/n44 ) );
  NAND3XL \DP_OP_725J1_134_142/U51  ( .A(\DP_OP_725J1_134_142/n42 ), .B(
        \DP_OP_725J1_134_142/n43 ), .C(\DP_OP_725J1_134_142/n44 ), .Y(
        \DP_OP_725J1_134_142/n224 ) );
  NAND2XL \DP_OP_725J1_134_142/U56  ( .A(N1677), .B(si_sel), .Y(
        \DP_OP_725J1_134_142/n45 ) );
  NAND2XL \DP_OP_725J1_134_142/U140  ( .A(\DP_OP_725J1_134_142/n262 ), .B(
        \DP_OP_725J1_134_142/I3 ), .Y(\DP_OP_725J1_134_142/n110 ) );
  NAND2XL \DP_OP_725J1_134_142/U142  ( .A(N752), .B(\DP_OP_725J1_134_142/I4 ), 
        .Y(\DP_OP_725J1_134_142/n112 ) );
  NAND2XL \DP_OP_725J1_134_142/U143  ( .A(n209), .B(\C169/Z_10 ), .Y(
        \DP_OP_725J1_134_142/n113 ) );
  NAND4XL \DP_OP_725J1_134_142/U139  ( .A(\DP_OP_725J1_134_142/n110 ), .B(
        \DP_OP_725J1_134_142/n111 ), .C(\DP_OP_725J1_134_142/n112 ), .D(
        \DP_OP_725J1_134_142/n113 ), .Y(\DP_OP_725J1_134_142/n243 ) );
  NAND2XL \DP_OP_725J1_134_142/U57  ( .A(\DP_OP_725J1_134_142/n243 ), .B(
        \DP_OP_725J1_134_142/I7 ), .Y(\DP_OP_725J1_134_142/n46 ) );
  NAND2XL \DP_OP_725J1_134_142/U58  ( .A(\DP_OP_725J1_134_142/I10 ), .B(
        \U3/RSOP_717/C2/Z_10 ), .Y(\DP_OP_725J1_134_142/n47 ) );
  NAND3XL \DP_OP_725J1_134_142/U55  ( .A(\DP_OP_725J1_134_142/n45 ), .B(
        \DP_OP_725J1_134_142/n46 ), .C(\DP_OP_725J1_134_142/n47 ), .Y(
        \DP_OP_725J1_134_142/n223 ) );
  NAND2XL \DP_OP_725J1_134_142/U60  ( .A(N1676), .B(si_sel), .Y(
        \DP_OP_725J1_134_142/n48 ) );
  NAND2XL \DP_OP_725J1_134_142/U145  ( .A(\DP_OP_725J1_134_142/n261 ), .B(
        \DP_OP_725J1_134_142/I3 ), .Y(\DP_OP_725J1_134_142/n114 ) );
  NAND2XL \DP_OP_725J1_134_142/U147  ( .A(N751), .B(\DP_OP_725J1_134_142/I4 ), 
        .Y(\DP_OP_725J1_134_142/n116 ) );
  NAND2XL \DP_OP_725J1_134_142/U148  ( .A(n209), .B(\C169/Z_9 ), .Y(
        \DP_OP_725J1_134_142/n117 ) );
  NAND4XL \DP_OP_725J1_134_142/U144  ( .A(\DP_OP_725J1_134_142/n114 ), .B(
        \DP_OP_725J1_134_142/n115 ), .C(\DP_OP_725J1_134_142/n116 ), .D(
        \DP_OP_725J1_134_142/n117 ), .Y(\DP_OP_725J1_134_142/n242 ) );
  NAND2XL \DP_OP_725J1_134_142/U61  ( .A(\DP_OP_725J1_134_142/n242 ), .B(
        \DP_OP_725J1_134_142/I7 ), .Y(\DP_OP_725J1_134_142/n49 ) );
  NAND2XL \DP_OP_725J1_134_142/U62  ( .A(\DP_OP_725J1_134_142/I10 ), .B(
        \U3/RSOP_717/C2/Z_9 ), .Y(\DP_OP_725J1_134_142/n50 ) );
  NAND3XL \DP_OP_725J1_134_142/U59  ( .A(\DP_OP_725J1_134_142/n48 ), .B(
        \DP_OP_725J1_134_142/n49 ), .C(\DP_OP_725J1_134_142/n50 ), .Y(
        \DP_OP_725J1_134_142/n222 ) );
  NAND2XL \DP_OP_725J1_134_142/U64  ( .A(N1675), .B(si_sel), .Y(
        \DP_OP_725J1_134_142/n51 ) );
  NAND2XL \DP_OP_725J1_134_142/U150  ( .A(\DP_OP_725J1_134_142/n260 ), .B(
        \DP_OP_725J1_134_142/I3 ), .Y(\DP_OP_725J1_134_142/n118 ) );
  NAND2XL \DP_OP_725J1_134_142/U152  ( .A(N750), .B(\DP_OP_725J1_134_142/I4 ), 
        .Y(\DP_OP_725J1_134_142/n120 ) );
  NAND2XL \DP_OP_725J1_134_142/U153  ( .A(n209), .B(\C169/Z_8 ), .Y(
        \DP_OP_725J1_134_142/n121 ) );
  NAND4XL \DP_OP_725J1_134_142/U149  ( .A(\DP_OP_725J1_134_142/n118 ), .B(
        \DP_OP_725J1_134_142/n119 ), .C(\DP_OP_725J1_134_142/n120 ), .D(
        \DP_OP_725J1_134_142/n121 ), .Y(\DP_OP_725J1_134_142/n241 ) );
  NAND2XL \DP_OP_725J1_134_142/U65  ( .A(\DP_OP_725J1_134_142/n241 ), .B(
        \DP_OP_725J1_134_142/I7 ), .Y(\DP_OP_725J1_134_142/n52 ) );
  NAND2XL \DP_OP_725J1_134_142/U66  ( .A(\DP_OP_725J1_134_142/I10 ), .B(
        \U3/RSOP_717/C2/Z_8 ), .Y(\DP_OP_725J1_134_142/n53 ) );
  NAND3XL \DP_OP_725J1_134_142/U63  ( .A(\DP_OP_725J1_134_142/n51 ), .B(
        \DP_OP_725J1_134_142/n52 ), .C(\DP_OP_725J1_134_142/n53 ), .Y(
        \DP_OP_725J1_134_142/n221 ) );
  NAND2XL \DP_OP_725J1_134_142/U68  ( .A(N1674), .B(si_sel), .Y(
        \DP_OP_725J1_134_142/n54 ) );
  XNOR2XL \DP_OP_725J1_134_142/U247  ( .A(\DP_OP_725J1_134_142/n202 ), .B(
        write_addr[9]), .Y(\DP_OP_725J1_134_142/n259 ) );
  NAND2XL \DP_OP_725J1_134_142/U156  ( .A(\DP_OP_725J1_134_142/n259 ), .B(
        \DP_OP_725J1_134_142/I3 ), .Y(\DP_OP_725J1_134_142/n123 ) );
  NAND3XL \DP_OP_725J1_134_142/U154  ( .A(\DP_OP_725J1_134_142/n122 ), .B(
        \DP_OP_725J1_134_142/n123 ), .C(\DP_OP_725J1_134_142/n124 ), .Y(
        \DP_OP_725J1_134_142/n240 ) );
  NAND2XL \DP_OP_725J1_134_142/U69  ( .A(\DP_OP_725J1_134_142/n240 ), .B(
        \DP_OP_725J1_134_142/I7 ), .Y(\DP_OP_725J1_134_142/n55 ) );
  NAND2XL \DP_OP_725J1_134_142/U70  ( .A(\DP_OP_725J1_134_142/I10 ), .B(
        \U3/RSOP_717/C2/Z_7 ), .Y(\DP_OP_725J1_134_142/n56 ) );
  NAND3XL \DP_OP_725J1_134_142/U67  ( .A(\DP_OP_725J1_134_142/n54 ), .B(
        \DP_OP_725J1_134_142/n55 ), .C(\DP_OP_725J1_134_142/n56 ), .Y(
        \DP_OP_725J1_134_142/n220 ) );
  NAND2XL \DP_OP_725J1_134_142/U72  ( .A(N1673), .B(si_sel), .Y(
        \DP_OP_725J1_134_142/n57 ) );
  NAND2XL \DP_OP_725J1_134_142/U159  ( .A(N627), .B(\DP_OP_725J1_134_142/I3 ), 
        .Y(\DP_OP_725J1_134_142/n125 ) );
  NAND3XL \DP_OP_725J1_134_142/U158  ( .A(\DP_OP_725J1_134_142/n126 ), .B(
        \DP_OP_725J1_134_142/n125 ), .C(\DP_OP_725J1_134_142/n127 ), .Y(
        \DP_OP_725J1_134_142/n239 ) );
  NAND2XL \DP_OP_725J1_134_142/U73  ( .A(\DP_OP_725J1_134_142/n239 ), .B(
        \DP_OP_725J1_134_142/I7 ), .Y(\DP_OP_725J1_134_142/n58 ) );
  NAND2XL \DP_OP_725J1_134_142/U74  ( .A(\DP_OP_725J1_134_142/I10 ), .B(
        \U3/RSOP_717/C2/Z_6 ), .Y(\DP_OP_725J1_134_142/n59 ) );
  NAND3XL \DP_OP_725J1_134_142/U71  ( .A(\DP_OP_725J1_134_142/n57 ), .B(
        \DP_OP_725J1_134_142/n58 ), .C(\DP_OP_725J1_134_142/n59 ), .Y(
        \DP_OP_725J1_134_142/n219 ) );
  NAND2XL \DP_OP_725J1_134_142/U76  ( .A(N1672), .B(si_sel), .Y(
        \DP_OP_725J1_134_142/n60 ) );
  NAND2XL \DP_OP_725J1_134_142/U163  ( .A(N626), .B(\DP_OP_725J1_134_142/I3 ), 
        .Y(\DP_OP_725J1_134_142/n128 ) );
  NAND3XL \DP_OP_725J1_134_142/U162  ( .A(\DP_OP_725J1_134_142/n129 ), .B(
        \DP_OP_725J1_134_142/n128 ), .C(\DP_OP_725J1_134_142/n130 ), .Y(
        \DP_OP_725J1_134_142/n238 ) );
  NAND2XL \DP_OP_725J1_134_142/U77  ( .A(\DP_OP_725J1_134_142/n238 ), .B(
        \DP_OP_725J1_134_142/I7 ), .Y(\DP_OP_725J1_134_142/n61 ) );
  NAND2XL \DP_OP_725J1_134_142/U78  ( .A(\DP_OP_725J1_134_142/I10 ), .B(
        \U3/RSOP_717/C2/Z_5 ), .Y(\DP_OP_725J1_134_142/n62 ) );
  NAND3XL \DP_OP_725J1_134_142/U75  ( .A(\DP_OP_725J1_134_142/n60 ), .B(
        \DP_OP_725J1_134_142/n61 ), .C(\DP_OP_725J1_134_142/n62 ), .Y(
        \DP_OP_725J1_134_142/n218 ) );
  NAND2XL \DP_OP_725J1_134_142/U80  ( .A(N1671), .B(si_sel), .Y(
        \DP_OP_725J1_134_142/n63 ) );
  NAND2XL \DP_OP_725J1_134_142/U167  ( .A(N625), .B(\DP_OP_725J1_134_142/I3 ), 
        .Y(\DP_OP_725J1_134_142/n131 ) );
  NAND3XL \DP_OP_725J1_134_142/U166  ( .A(\DP_OP_725J1_134_142/n132 ), .B(
        \DP_OP_725J1_134_142/n131 ), .C(\DP_OP_725J1_134_142/n133 ), .Y(
        \DP_OP_725J1_134_142/n237 ) );
  NAND2XL \DP_OP_725J1_134_142/U81  ( .A(\DP_OP_725J1_134_142/n237 ), .B(
        \DP_OP_725J1_134_142/I7 ), .Y(\DP_OP_725J1_134_142/n64 ) );
  NAND2XL \DP_OP_725J1_134_142/U82  ( .A(\DP_OP_725J1_134_142/I10 ), .B(
        \U3/RSOP_717/C2/Z_4 ), .Y(\DP_OP_725J1_134_142/n65 ) );
  NAND3XL \DP_OP_725J1_134_142/U79  ( .A(\DP_OP_725J1_134_142/n63 ), .B(
        \DP_OP_725J1_134_142/n64 ), .C(\DP_OP_725J1_134_142/n65 ), .Y(
        \DP_OP_725J1_134_142/n217 ) );
  NAND2XL \DP_OP_725J1_134_142/U84  ( .A(N1670), .B(si_sel), .Y(
        \DP_OP_725J1_134_142/n66 ) );
  NAND2XL \DP_OP_725J1_134_142/U171  ( .A(N624), .B(\DP_OP_725J1_134_142/I3 ), 
        .Y(\DP_OP_725J1_134_142/n134 ) );
  NAND3XL \DP_OP_725J1_134_142/U170  ( .A(\DP_OP_725J1_134_142/n135 ), .B(
        \DP_OP_725J1_134_142/n134 ), .C(\DP_OP_725J1_134_142/n136 ), .Y(
        \DP_OP_725J1_134_142/n236 ) );
  NAND2XL \DP_OP_725J1_134_142/U85  ( .A(\DP_OP_725J1_134_142/n236 ), .B(
        \DP_OP_725J1_134_142/I7 ), .Y(\DP_OP_725J1_134_142/n67 ) );
  NAND2XL \DP_OP_725J1_134_142/U86  ( .A(\DP_OP_725J1_134_142/I10 ), .B(
        \U3/RSOP_717/C2/Z_3 ), .Y(\DP_OP_725J1_134_142/n68 ) );
  NAND3XL \DP_OP_725J1_134_142/U83  ( .A(\DP_OP_725J1_134_142/n66 ), .B(
        \DP_OP_725J1_134_142/n67 ), .C(\DP_OP_725J1_134_142/n68 ), .Y(
        \DP_OP_725J1_134_142/n216 ) );
  NAND2XL \DP_OP_725J1_134_142/U88  ( .A(N1669), .B(si_sel), .Y(
        \DP_OP_725J1_134_142/n69 ) );
  NAND2XL \DP_OP_725J1_134_142/U175  ( .A(N623), .B(\DP_OP_725J1_134_142/I3 ), 
        .Y(\DP_OP_725J1_134_142/n137 ) );
  NAND3XL \DP_OP_725J1_134_142/U174  ( .A(\DP_OP_725J1_134_142/n138 ), .B(
        \DP_OP_725J1_134_142/n137 ), .C(n107), .Y(\DP_OP_725J1_134_142/n235 )
         );
  NAND2XL \DP_OP_725J1_134_142/U89  ( .A(\DP_OP_725J1_134_142/n235 ), .B(
        \DP_OP_725J1_134_142/I7 ), .Y(\DP_OP_725J1_134_142/n70 ) );
  NAND2XL \DP_OP_725J1_134_142/U90  ( .A(\DP_OP_725J1_134_142/I10 ), .B(
        \U3/RSOP_717/C2/Z_2 ), .Y(\DP_OP_725J1_134_142/n71 ) );
  NAND3XL \DP_OP_725J1_134_142/U87  ( .A(\DP_OP_725J1_134_142/n69 ), .B(
        \DP_OP_725J1_134_142/n70 ), .C(\DP_OP_725J1_134_142/n71 ), .Y(
        \DP_OP_725J1_134_142/n215 ) );
  NAND2XL \DP_OP_725J1_134_142/U182  ( .A(\DP_OP_725J1_134_142/n143 ), .B(
        \DP_OP_725J1_134_142/n144 ), .Y(\DP_OP_725J1_134_142/n233 ) );
  NAND2XL \DP_OP_725J1_134_142/U96  ( .A(\DP_OP_725J1_134_142/n233 ), .B(
        \DP_OP_725J1_134_142/I7 ), .Y(\DP_OP_725J1_134_142/n75 ) );
  NAND2XL \DP_OP_725J1_134_142/U97  ( .A(N1667), .B(si_sel), .Y(
        \DP_OP_725J1_134_142/n76 ) );
  NAND2XL \DP_OP_725J1_134_142/U98  ( .A(\DP_OP_725J1_134_142/I10 ), .B(
        \U3/RSOP_717/C2/Z_0 ), .Y(\DP_OP_725J1_134_142/n77 ) );
  NAND3XL \DP_OP_725J1_134_142/U95  ( .A(\DP_OP_725J1_134_142/n75 ), .B(
        \DP_OP_725J1_134_142/n76 ), .C(\DP_OP_725J1_134_142/n77 ), .Y(
        \DP_OP_725J1_134_142/n213 ) );
  NAND2XL \DP_OP_725J1_134_142/U92  ( .A(N1668), .B(si_sel), .Y(
        \DP_OP_725J1_134_142/n72 ) );
  NAND2XL \DP_OP_725J1_134_142/U179  ( .A(N622), .B(\DP_OP_725J1_134_142/I3 ), 
        .Y(\DP_OP_725J1_134_142/n140 ) );
  NAND3XL \DP_OP_725J1_134_142/U178  ( .A(\DP_OP_725J1_134_142/n141 ), .B(
        \DP_OP_725J1_134_142/n140 ), .C(\DP_OP_725J1_134_142/n142 ), .Y(
        \DP_OP_725J1_134_142/n234 ) );
  NAND2XL \DP_OP_725J1_134_142/U93  ( .A(\DP_OP_725J1_134_142/n234 ), .B(
        \DP_OP_725J1_134_142/I7 ), .Y(\DP_OP_725J1_134_142/n73 ) );
  NAND2XL \DP_OP_725J1_134_142/U94  ( .A(\DP_OP_725J1_134_142/I10 ), .B(
        \U3/RSOP_717/C2/Z_1 ), .Y(\DP_OP_725J1_134_142/n74 ) );
  NAND3XL \DP_OP_725J1_134_142/U91  ( .A(\DP_OP_725J1_134_142/n72 ), .B(
        \DP_OP_725J1_134_142/n73 ), .C(\DP_OP_725J1_134_142/n74 ), .Y(
        \DP_OP_725J1_134_142/n214 ) );
  XOR2XL \DP_OP_725J1_134_142/U186  ( .A(write_addr[19]), .B(fb_addr[19]), .Y(
        \DP_OP_725J1_134_142/n145 ) );
  XOR2XL \DP_OP_725J1_134_142/U2  ( .A(\DP_OP_725J1_134_142/n232 ), .B(
        \C1/Z_19 ), .Y(\DP_OP_725J1_134_142/n1 ) );
  XOR2XL \DP_OP_725J1_134_142/U1  ( .A(\DP_OP_725J1_134_142/n2 ), .B(
        \DP_OP_725J1_134_142/n1 ), .Y(\C168/DATA3_19 ) );
  AND2XL \DP_OP_280J1_126_7605/U12  ( .A(\C1/Z_0 ), .B(n85), .Y(
        \DP_OP_280J1_126_7605/n16 ) );
  AND2XL \DP_OP_280J1_126_7605/U7  ( .A(\DP_OP_280J1_126_7605/n27 ), .B(n85), 
        .Y(\DP_OP_280J1_126_7605/n21 ) );
  DFFRX4 \work_cntr_reg[4]  ( .D(next_work_cntr[4]), .CK(clk), .RN(n43), .Q(
        work_cntr[4]), .QN(n164) );
  DFFRX2 \work_cntr_reg[5]  ( .D(next_work_cntr[5]), .CK(clk), .RN(n43), .Q(
        work_cntr[5]), .QN(n197) );
  DFFRX4 \work_cntr_reg[2]  ( .D(next_work_cntr[2]), .CK(clk), .RN(n43), .Q(
        N2283), .QN(n199) );
  DFFRX2 \work_cntr_reg[17]  ( .D(next_work_cntr[17]), .CK(clk), .RN(n43), .Q(
        work_cntr[17]), .QN(n182) );
  DFFRX2 \work_cntr_reg[15]  ( .D(next_work_cntr[15]), .CK(clk), .RN(n43), .Q(
        work_cntr[15]), .QN(n188) );
  DFFRX2 \write_cntr_reg/q_reg[10]  ( .D(n537), .CK(clk), .RN(n43), .Q(
        write_cntr[10]), .QN(n204) );
  DFFRX2 \work_cntr_reg[9]  ( .D(next_work_cntr[9]), .CK(clk), .RN(n43), .Q(
        work_cntr[9]), .QN(n187) );
  DFFRX2 \write_addr_reg/q_reg[9]  ( .D(n492), .CK(clk), .RN(n43), .Q(
        write_addr[9]), .QN(n233) );
  DFFRXL \write_addr_reg/q_reg[12]  ( .D(n489), .CK(clk), .RN(n43), .Q(
        write_addr[12]), .QN(n236) );
  DFFRX4 \write_addr_reg/q_reg[16]  ( .D(n485), .CK(clk), .RN(n43), .Q(
        write_addr[16]), .QN(n239) );
  ADDHX1 \DP_OP_725J1_134_142/U221  ( .A(write_addr[16]), .B(
        \DP_OP_725J1_134_142/n178 ), .CO(\DP_OP_725J1_134_142/n177 ), .S(N635)
         );
  ADDHX1 \DP_OP_725J1_134_142/U209  ( .A(write_addr[16]), .B(
        \DP_OP_725J1_134_142/n168 ), .CO(\DP_OP_725J1_134_142/n167 ), .S(N756)
         );
  DFFRX4 \read_cntr_reg/q_reg[0]  ( .D(n521), .CK(clk), .RN(n43), .Q(
        read_cntr[0]), .QN(n171) );
  DFFRX2 \write_cntr_reg/q_reg[5]  ( .D(n541), .CK(clk), .RN(n43), .Q(
        write_cntr[5]), .QN(n198) );
  DFFRX2 \write_cntr_reg/q_reg[8]  ( .D(n545), .CK(clk), .RN(n43), .Q(
        write_cntr[8]), .QN(n195) );
  DFFRX2 \work_cntr_reg[0]  ( .D(next_work_cntr[0]), .CK(clk), .RN(n43), .Q(
        N205), .QN(n146) );
  DFFRX2 \write_cntr_reg/q_reg[7]  ( .D(n539), .CK(clk), .RN(n43), .Q(
        write_cntr[7]), .QN(n196) );
  DFFRX4 \work_cntr_reg[13]  ( .D(next_work_cntr[13]), .CK(clk), .RN(n43), .Q(
        work_cntr[13]), .QN(n184) );
  DFFRX4 \write_addr_reg/q_reg[18]  ( .D(n483), .CK(clk), .RN(n43), .Q(
        write_addr[18]), .QN(n246) );
  ADDHX1 \DP_OP_725J1_134_142/U219  ( .A(write_addr[18]), .B(
        \DP_OP_725J1_134_142/n176 ), .CO(\DP_OP_725J1_134_142/n175 ), .S(N637)
         );
  ADDHX1 \DP_OP_725J1_134_142/U207  ( .A(write_addr[18]), .B(
        \DP_OP_725J1_134_142/n166 ), .CO(\DP_OP_725J1_134_142/n165 ), .S(N758)
         );
  DFFRX2 \write_addr_reg/q_reg[11]  ( .D(n490), .CK(clk), .RN(n802), .Q(
        write_addr[11]), .QN(n153) );
  DFFRX2 \work_cntr_reg[10]  ( .D(next_work_cntr[10]), .CK(clk), .RN(n43), .Q(
        work_cntr[10]), .QN(n160) );
  DFFRX2 \work_cntr_reg[19]  ( .D(next_work_cntr[19]), .CK(clk), .RN(n802), 
        .Q(work_cntr[19]), .QN(n152) );
  DFFRX2 \write_addr_reg/q_reg[5]  ( .D(n525), .CK(clk), .RN(n802), .Q(N746), 
        .QN(n213) );
  DFFRX2 \write_addr_reg/q_reg[8]  ( .D(n493), .CK(clk), .RN(n802), .Q(
        write_addr[8]), .QN(n207) );
  DFFRX2 \work_cntr_reg[16]  ( .D(next_work_cntr[16]), .CK(clk), .RN(n43), .Q(
        work_cntr[16]), .QN(n181) );
  DFFRX2 \write_addr_reg/q_reg[15]  ( .D(n486), .CK(clk), .RN(n802), .Q(
        write_addr[15]), .QN(n234) );
  ADDHX1 \DP_OP_725J1_134_142/U222  ( .A(write_addr[15]), .B(
        \DP_OP_725J1_134_142/n179 ), .CO(\DP_OP_725J1_134_142/n178 ), .S(N634)
         );
  ADDHX1 \DP_OP_725J1_134_142/U210  ( .A(write_addr[15]), .B(
        \DP_OP_725J1_134_142/n169 ), .CO(\DP_OP_725J1_134_142/n168 ), .S(N755)
         );
  DFFRX4 \write_addr_reg/q_reg[10]  ( .D(n491), .CK(clk), .RN(n43), .Q(
        write_addr[10]), .QN(n169) );
  ADDHX1 \DP_OP_725J1_134_142/U227  ( .A(write_addr[10]), .B(
        \DP_OP_725J1_134_142/n184 ), .CO(\DP_OP_725J1_134_142/n183 ), .S(N629)
         );
  ADDHX1 \DP_OP_725J1_134_142/U215  ( .A(write_addr[10]), .B(write_addr[9]), 
        .CO(\DP_OP_725J1_134_142/n173 ), .S(N750) );
  DFFSX2 \state_reg[0]  ( .D(n781), .CK(clk), .SN(n43), .Q(n163), .QN(state[0]) );
  DFFRX2 \write_addr_reg/q_reg[7]  ( .D(n523), .CK(clk), .RN(n43), .Q(N748), 
        .QN(n168) );
  ADDHX1 \DP_OP_725J1_134_142/U249  ( .A(N748), .B(\DP_OP_725J1_134_142/n203 ), 
        .CO(\DP_OP_725J1_134_142/n202 ), .S(N627) );
  DFFRX2 \write_addr_reg/q_reg[1]  ( .D(n529), .CK(clk), .RN(n43), .Q(N742), 
        .QN(n173) );
  DFFRX2 \work_cntr_reg[18]  ( .D(next_work_cntr[18]), .CK(clk), .RN(n43), .Q(
        work_cntr[18]), .QN(n161) );
  DFFRX4 \work_cntr_reg[3]  ( .D(next_work_cntr[3]), .CK(clk), .RN(n43), .Q(
        N2284), .QN(n162) );
  DFFRX2 \write_addr_reg/q_reg[2]  ( .D(n528), .CK(clk), .RN(n43), .Q(N743), 
        .QN(n137) );
  ADDHX1 \DP_OP_725J1_134_142/U234  ( .A(N743), .B(N742), .CO(
        \DP_OP_725J1_134_142/n190 ), .S(N622) );
  DFFRX2 \write_addr_reg/q_reg[3]  ( .D(n527), .CK(clk), .RN(n802), .Q(N744), 
        .QN(n211) );
  ADDHX1 \DP_OP_725J1_134_142/U253  ( .A(N744), .B(\DP_OP_725J1_134_142/n190 ), 
        .CO(\DP_OP_725J1_134_142/n206 ), .S(N623) );
  ADDHX1 \DP_OP_725J1_134_142/U231  ( .A(N746), .B(\DP_OP_725J1_134_142/n205 ), 
        .CO(\DP_OP_725J1_134_142/n187 ), .S(N625) );
  ADDHX1 \DP_OP_725J1_134_142/U250  ( .A(N747), .B(\DP_OP_725J1_134_142/n187 ), 
        .CO(\DP_OP_725J1_134_142/n203 ), .S(N626) );
  ADDHX1 \DP_OP_725J1_134_142/U252  ( .A(N745), .B(\DP_OP_725J1_134_142/n206 ), 
        .CO(\DP_OP_725J1_134_142/n205 ), .S(N624) );
  DFFRX2 \write_addr_reg/q_reg[17]  ( .D(n484), .CK(clk), .RN(n43), .Q(
        write_addr[17]), .QN(n154) );
  DFFRX2 \write_addr_reg/q_reg[19]  ( .D(n482), .CK(clk), .RN(n802), .Q(
        write_addr[19]), .QN(n208) );
  DFFRX2 \write_cntr_reg/q_reg[13]  ( .D(n534), .CK(clk), .RN(n43), .Q(
        write_cntr[13]), .QN(n202) );
  ADDHX1 \DP_OP_725J1_134_142/U205  ( .A(fb_addr[0]), .B(
        \next_write_addr_w[0] ), .CO(\DP_OP_725J1_134_142/n164 ), .S(N1667) );
  ADDHX1 \DP_OP_725J1_134_142/U213  ( .A(n102), .B(\DP_OP_725J1_134_142/n172 ), 
        .CO(\DP_OP_725J1_134_142/n171 ), .S(N752) );
  ADDHX1 \DP_OP_725J1_134_142/U214  ( .A(write_addr[11]), .B(
        \DP_OP_725J1_134_142/n173 ), .CO(\DP_OP_725J1_134_142/n172 ), .S(N751)
         );
  ADDHX1 \DP_OP_725J1_134_142/U212  ( .A(n89), .B(\DP_OP_725J1_134_142/n171 ), 
        .CO(\DP_OP_725J1_134_142/n170 ), .S(N753) );
  DFFRX2 \write_addr_reg/q_reg[6]  ( .D(n524), .CK(clk), .RN(n43), .Q(N747), 
        .QN(n136) );
  DFFRX4 \work_cntr_reg[11]  ( .D(next_work_cntr[11]), .CK(clk), .RN(n43), .Q(
        work_cntr[11]), .QN(n180) );
  DFFRX2 \write_addr_reg/q_reg[4]  ( .D(n526), .CK(clk), .RN(n43), .Q(N745), 
        .QN(n167) );
  ADDHX1 \DP_OP_725J1_134_142/U225  ( .A(n102), .B(\DP_OP_725J1_134_142/n182 ), 
        .CO(\DP_OP_725J1_134_142/n181 ), .S(N631) );
  ADDHX1 \DP_OP_725J1_134_142/U224  ( .A(n89), .B(\DP_OP_725J1_134_142/n181 ), 
        .CO(\DP_OP_725J1_134_142/n180 ), .S(N632) );
  ADDHX1 \DP_OP_725J1_134_142/U220  ( .A(write_addr[17]), .B(
        \DP_OP_725J1_134_142/n177 ), .CO(\DP_OP_725J1_134_142/n176 ), .S(N636)
         );
  ADDHX1 \DP_OP_725J1_134_142/U218  ( .A(write_addr[19]), .B(
        \DP_OP_725J1_134_142/n175 ), .CO(N639), .S(N638) );
  ADDHX1 \DP_OP_725J1_134_142/U226  ( .A(write_addr[11]), .B(
        \DP_OP_725J1_134_142/n183 ), .CO(\DP_OP_725J1_134_142/n182 ), .S(N630)
         );
  ADDHX1 \DP_OP_725J1_134_142/U228  ( .A(write_addr[9]), .B(
        \DP_OP_725J1_134_142/n202 ), .CO(\DP_OP_725J1_134_142/n184 ), .S(N628)
         );
  ADDHX1 \DP_OP_725J1_134_142/U211  ( .A(n88), .B(\DP_OP_725J1_134_142/n170 ), 
        .CO(\DP_OP_725J1_134_142/n169 ), .S(N754) );
  ADDHX1 \DP_OP_725J1_134_142/U208  ( .A(write_addr[17]), .B(
        \DP_OP_725J1_134_142/n167 ), .CO(\DP_OP_725J1_134_142/n166 ), .S(N757)
         );
  ADDHX1 \DP_OP_725J1_134_142/U206  ( .A(write_addr[19]), .B(
        \DP_OP_725J1_134_142/n165 ), .CO(N760), .S(N759) );
  DFFRX4 \work_cntr_reg[1]  ( .D(next_work_cntr[1]), .CK(clk), .RN(n43), .Q(
        N2282), .QN(n165) );
  DFFRX2 \write_cntr_reg/q_reg[11]  ( .D(n536), .CK(clk), .RN(n43), .Q(
        write_cntr[11]), .QN(n189) );
  DFFRX2 \write_cntr_reg/q_reg[4]  ( .D(n546), .CK(clk), .RN(n43), .Q(
        write_cntr[4]), .QN(n166) );
  DFFRX2 \work_cntr_reg[12]  ( .D(next_work_cntr[12]), .CK(clk), .RN(n802), 
        .Q(work_cntr[12]), .QN(n2548) );
  DFFRX2 \work_cntr_reg[6]  ( .D(next_work_cntr[6]), .CK(clk), .RN(n802), .Q(
        work_cntr[6]), .QN(n2600) );
  DFFRX1 en_si_reg ( .D(n2931), .CK(clk), .RN(n43), .QN(en_si) );
  DFFRX1 \global_cntr_reg[0]  ( .D(n183), .CK(clk), .RN(n802), .Q(
        global_cntr[0]), .QN(n183) );
  DFFRX1 \global_cntr_reg[1]  ( .D(\next_glb_cntr[1] ), .CK(clk), .RN(n43), 
        .Q(global_cntr[1]), .QN(n155) );
  DFFRX1 \global_cntr_reg[2]  ( .D(n797), .CK(clk), .RN(n802), .Q(
        global_cntr[2]), .QN(n150) );
  DFFRX1 \global_cntr_reg[3]  ( .D(n795), .CK(clk), .RN(n802), .Q(
        global_cntr[3]), .QN(n156) );
  DFFRX1 \global_cntr_reg[4]  ( .D(n794), .CK(clk), .RN(n802), .Q(
        global_cntr[4]), .QN(n138) );
  DFFRX1 \global_cntr_reg[5]  ( .D(n793), .CK(clk), .RN(n802), .Q(
        global_cntr[5]), .QN(n157) );
  DFFRX1 \global_cntr_reg[6]  ( .D(n792), .CK(clk), .RN(n802), .Q(
        global_cntr[6]), .QN(n139) );
  DFFRX1 \global_cntr_reg[7]  ( .D(n791), .CK(clk), .RN(n802), .Q(
        global_cntr[7]), .QN(n158) );
  DFFRX1 \global_cntr_reg[8]  ( .D(n790), .CK(clk), .RN(n802), .Q(
        global_cntr[8]), .QN(n142) );
  DFFRX1 \global_cntr_reg[9]  ( .D(n789), .CK(clk), .RN(n802), .Q(
        global_cntr[9]), .QN(n147) );
  DFFRX1 \global_cntr_reg[11]  ( .D(n787), .CK(clk), .RN(n802), .Q(
        global_cntr[11]), .QN(n141) );
  DFFRX1 \global_cntr_reg[10]  ( .D(n788), .CK(clk), .RN(n802), .Q(
        global_cntr[10]), .QN(n159) );
  DFFRX1 \global_cntr_reg[12]  ( .D(n801), .CK(clk), .RN(n802), .Q(
        global_cntr[12]), .QN(n174) );
  DFFRX1 \global_cntr_reg[13]  ( .D(n800), .CK(clk), .RN(n802), .Q(
        global_cntr[13]), .QN(n143) );
  DFFRX1 \global_cntr_reg[15]  ( .D(n786), .CK(clk), .RN(n802), .Q(
        global_cntr[15]), .QN(n144) );
  DFFRX1 \global_cntr_reg[14]  ( .D(n799), .CK(clk), .RN(n802), .Q(
        global_cntr[14]), .QN(n145) );
  DFFRX1 \global_cntr_reg[16]  ( .D(n785), .CK(clk), .RN(n802), .Q(
        global_cntr[16]), .QN(n140) );
  DFFRX1 \global_cntr_reg[19]  ( .D(n782), .CK(clk), .RN(n802), .Q(
        global_cntr[19]), .QN(n176) );
  DFFRX1 \global_cntr_reg[18]  ( .D(n783), .CK(clk), .RN(n802), .Q(
        global_cntr[18]), .QN(n149) );
  DFFRX1 \global_cntr_reg[17]  ( .D(n784), .CK(clk), .RN(n802), .Q(
        global_cntr[17]), .QN(n148) );
  DFFRX1 \state_reg[1]  ( .D(next_state[1]), .CK(clk), .RN(n802), .Q(n185), 
        .QN(n32) );
  DFFRX1 \state_reg[2]  ( .D(next_state[2]), .CK(clk), .RN(n802), .Q(state[2]), 
        .QN(n190) );
  DFFRX1 \work_cntr_reg[7]  ( .D(next_work_cntr[7]), .CK(clk), .RN(n802), .Q(
        work_cntr[7]), .QN(n194) );
  DFFRX1 \curr_photo_reg[1]  ( .D(next_photo[1]), .CK(clk), .RN(n802), .Q(
        curr_photo[1]), .QN(n243) );
  DFFRX1 \curr_photo_reg[0]  ( .D(next_photo[0]), .CK(clk), .RN(n802), .Q(
        curr_photo[0]), .QN(n244) );
  DFFRX1 \write_cntr_reg/q_reg[6]  ( .D(n540), .CK(clk), .RN(n802), .Q(
        write_cntr[6]), .QN(n191) );
  DFFRX1 \write_cntr_reg/q_reg[3]  ( .D(n542), .CK(clk), .RN(n802), .Q(
        write_cntr[3]), .QN(n200) );
  DFFRX1 \write_cntr_reg/q_reg[0]  ( .D(n543), .CK(clk), .RN(n802), .Q(
        write_cntr[0]), .QN(n203) );
  DFFRX1 \write_cntr_reg/q_reg[14]  ( .D(n533), .CK(clk), .RN(n802), .Q(
        write_cntr[14]), .QN(n205) );
  DFFRX1 \write_cntr_reg/q_reg[9]  ( .D(n538), .CK(clk), .RN(n802), .Q(
        write_cntr[9]), .QN(n192) );
  DFFRX1 \write_addr_reg/q_reg[14]  ( .D(n487), .CK(clk), .RN(n802), .Q(
        write_addr[14]), .QN(n235) );
  DFFRX1 \write_addr_reg/q_reg[0]  ( .D(n530), .CK(clk), .RN(n802), .Q(
        \next_write_addr_w[0] ), .QN(n212) );
  DFFRX1 \write_cntr_reg/q_reg[1]  ( .D(n548), .CK(clk), .RN(n802), .Q(
        write_cntr[1]), .QN(n201) );
  DFFRX1 \write_addr_reg/q_reg[13]  ( .D(n488), .CK(clk), .RN(n802), .Q(
        write_addr[13]), .QN(n206) );
  DFFRX1 \read_cntr_reg/q_reg[1]  ( .D(n520), .CK(clk), .RN(n802), .Q(
        read_cntr[1]), .QN(n172) );
  DFFRX1 \cr_read_cntr_reg/q_reg[1]  ( .D(n501), .CK(clk), .RN(n802), .Q(N1454), .QN(n245) );
  DFFRX1 \cr_read_cntr_reg/q_reg[3]  ( .D(n499), .CK(clk), .RN(n802), .Q(
        cr_read_cntr[3]), .QN(n240) );
  DFFRX1 \cr_read_cntr_reg/q_reg[4]  ( .D(n498), .CK(clk), .RN(n802), .Q(
        cr_read_cntr[4]), .QN(n241) );
  DFFRX1 \cr_read_cntr_reg/q_reg[5]  ( .D(n497), .CK(clk), .RN(n802), .Q(
        cr_read_cntr[5]), .QN(n238) );
  DFFRX1 \cr_read_cntr_reg/q_reg[6]  ( .D(n496), .CK(clk), .RN(n802), .Q(
        cr_read_cntr[6]), .QN(n242) );
  DFFRX1 \work_cntr_reg[14]  ( .D(next_work_cntr[14]), .CK(clk), .RN(n43), .Q(
        work_cntr[14]) );
  DFFRX1 \write_cntr_reg/q_reg[2]  ( .D(n547), .CK(clk), .RN(n43), .Q(
        write_cntr[2]), .QN(n3) );
  DFFRX1 \cr_read_cntr_reg/q_reg[0]  ( .D(n502), .CK(clk), .RN(n43), .Q(N1453), 
        .QN(n6) );
  DFFRX1 \cr_read_cntr_reg/q_reg[2]  ( .D(n500), .CK(clk), .RN(n43), .Q(N1455), 
        .QN(n9) );
  DFFRX2 \write_cntr_reg/q_reg[12]  ( .D(n535), .CK(clk), .RN(n802), .Q(
        write_cntr[12]), .QN(n2144) );
  DFFRX2 \work_cntr_reg[8]  ( .D(next_work_cntr[8]), .CK(clk), .RN(n43), .Q(
        work_cntr[8]), .QN(n193) );
  NAND2X1 U3 ( .A(n1998), .B(n1997), .Y(n2005) );
  OR2X1 U4 ( .A(n164), .B(n2149), .Y(n1) );
  OR2X1 U5 ( .A(n974), .B(n973), .Y(n2) );
  AOI211X1 U6 ( .A0(n2018), .A1(n2017), .B0(n2016), .C0(n2015), .Y(n2028) );
  NAND2X1 U7 ( .A(n2833), .B(n2832), .Y(n2867) );
  AOI2BB1X1 U8 ( .A0N(n161), .A1N(n1726), .B0(n1731), .Y(n1735) );
  OAI2BB1X1 U9 ( .A0N(n197), .A1N(n1), .B0(n1045), .Y(n2450) );
  OAI21XL U10 ( .A0(n2322), .A1(n163), .B0(n840), .Y(n178) );
  CLKINVX1 U11 ( .A(curr_photo_size[0]), .Y(n2923) );
  NAND2BX1 U12 ( .AN(state[0]), .B(en_so), .Y(n2122) );
  OAI2BB1X1 U13 ( .A0N(n2), .A1N(n3), .B0(n975), .Y(n2133) );
  NOR2X1 U14 ( .A(n144), .B(n272), .Y(n273) );
  NOR2X1 U15 ( .A(n263), .B(n138), .Y(n264) );
  OAI2BB2XL U16 ( .B0(n1377), .B1(n1376), .A0N(n1377), .A1N(n1376), .Y(n4) );
  CLKBUFX3 U17 ( .A(n2945), .Y(n42) );
  BUFX4 U18 ( .A(n178), .Y(n41) );
  NOR2X1 U19 ( .A(n2100), .B(n2969), .Y(expand_sel[2]) );
  OR2X1 U20 ( .A(n6), .B(n2969), .Y(n5) );
  OR2X1 U21 ( .A(n245), .B(n2969), .Y(n7) );
  OR2X1 U22 ( .A(n9), .B(n2969), .Y(n8) );
  OR2X1 U23 ( .A(n11), .B(n2969), .Y(n10) );
  XNOR2X1 U24 ( .A(\DP_OP_280J1_126_7605/n1 ), .B(\DP_OP_280J1_126_7605/n21 ), 
        .Y(n11) );
  CLKAND2X3 U25 ( .A(n621), .B(n620), .Y(n718) );
  NOR2X2 U26 ( .A(n2122), .B(n2923), .Y(n669) );
  NAND3X1 U27 ( .A(n2500), .B(n1254), .C(n2600), .Y(n1226) );
  NOR2X1 U28 ( .A(n2715), .B(n2713), .Y(n12) );
  AOI2BB2X1 U29 ( .B0(n2714), .B1(n12), .A0N(n2714), .A1N(n12), .Y(n2737) );
  OAI2BB1X1 U30 ( .A0N(n1903), .A1N(n1902), .B0(n1901), .Y(n1950) );
  AO21X1 U31 ( .A0(\DP_OP_280J1_126_7605/n25 ), .A1(n85), .B0(
        \DP_OP_280J1_126_7605/I2 ), .Y(n13) );
  AND2X1 U32 ( .A(\DP_OP_280J1_126_7605/n3 ), .B(n13), .Y(
        \DP_OP_280J1_126_7605/n2 ) );
  AOI2BB2X1 U33 ( .B0(\DP_OP_280J1_126_7605/n3 ), .B1(n13), .A0N(
        \DP_OP_280J1_126_7605/n3 ), .A1N(n13), .Y(N1459) );
  NOR4X1 U34 ( .A(n2741), .B(n48), .C(n2720), .D(n2716), .Y(n14) );
  NAND3X1 U35 ( .A(n2735), .B(n2733), .C(n14), .Y(n2739) );
  OAI2BB1X1 U36 ( .A0N(n1905), .A1N(n1914), .B0(n1915), .Y(n1949) );
  AO21X1 U37 ( .A0(\DP_OP_280J1_126_7605/n26 ), .A1(n85), .B0(
        \DP_OP_280J1_126_7605/I2 ), .Y(n15) );
  AND2X1 U38 ( .A(\DP_OP_280J1_126_7605/n2 ), .B(n15), .Y(
        \DP_OP_280J1_126_7605/n1 ) );
  AOI2BB2X1 U39 ( .B0(\DP_OP_280J1_126_7605/n2 ), .B1(n15), .A0N(
        \DP_OP_280J1_126_7605/n2 ), .A1N(n15), .Y(N1460) );
  NOR2X1 U40 ( .A(n2729), .B(n2736), .Y(n16) );
  AOI2BB2X1 U41 ( .B0(n77), .B1(n16), .A0N(n77), .A1N(n16), .Y(n2753) );
  OAI21XL U42 ( .A0(n2829), .A1(n2775), .B0(n2774), .Y(n17) );
  XNOR2X1 U43 ( .A(n17), .B(n2776), .Y(n2802) );
  NAND2X1 U44 ( .A(n859), .B(next_cr_x[6]), .Y(n18) );
  XNOR2X1 U45 ( .A(n18), .B(n869), .Y(n1050) );
  NAND3BX1 U46 ( .AN(n1868), .B(n1710), .C(read_cntr[1]), .Y(n506) );
  OAI2BB1X1 U47 ( .A0N(n1891), .A1N(n1888), .B0(n1889), .Y(n1951) );
  OAI2BB1X1 U48 ( .A0N(n1929), .A1N(n1927), .B0(n1919), .Y(n2131) );
  OAI21XL U49 ( .A0(n78), .A1(n2777), .B0(n2757), .Y(n19) );
  XNOR2X1 U50 ( .A(n19), .B(n2758), .Y(n2794) );
  NAND3X1 U51 ( .A(n2829), .B(n2828), .C(n2827), .Y(n20) );
  AOI2BB2X1 U52 ( .B0(n2830), .B1(n20), .A0N(n2830), .A1N(n20), .Y(n2857) );
  AOI31X1 U53 ( .A0(n869), .A1(next_cr_x[6]), .A2(n859), .B0(n867), .Y(n1060)
         );
  NAND2BX1 U54 ( .AN(curr_time[1]), .B(n428), .Y(n429) );
  OAI2BB1X1 U55 ( .A0N(n981), .A1N(n984), .B0(n977), .Y(n1375) );
  AO21X1 U56 ( .A0(n2959), .A1(n146), .B0(n1864), .Y(n21) );
  NAND2X1 U57 ( .A(n2644), .B(n199), .Y(n22) );
  NAND3X1 U58 ( .A(n619), .B(n21), .C(n22), .Y(n623) );
  NOR2BX1 U59 ( .AN(n669), .B(curr_photo_size[1]), .Y(n766) );
  NOR2X1 U60 ( .A(n2129), .B(n2128), .Y(n23) );
  NAND2X1 U61 ( .A(n381), .B(n23), .Y(n465) );
  NOR2X1 U62 ( .A(n359), .B(N1455), .Y(n24) );
  AOI211X1 U63 ( .A0(n359), .A1(N1455), .B0(n41), .C0(n24), .Y(n500) );
  XNOR2X1 U64 ( .A(n2703), .B(n2702), .Y(n48) );
  OAI2BB1X1 U65 ( .A0N(n113), .A1N(n2020), .B0(n2005), .Y(n2017) );
  NOR2X1 U66 ( .A(n2732), .B(n2730), .Y(n25) );
  AOI2BB2X1 U67 ( .B0(n2731), .B1(n25), .A0N(n2731), .A1N(n25), .Y(n2764) );
  AOI2BB2X1 U68 ( .B0(n2813), .B1(n2812), .A0N(n2813), .A1N(n2812), .Y(n26) );
  XNOR2X1 U69 ( .A(n26), .B(n2814), .Y(n2845) );
  CLKINVX1 U70 ( .A(n1336), .Y(n27) );
  AOI32X1 U71 ( .A0(n1334), .A1(n27), .A2(n1333), .B0(n1336), .B1(n1335), .Y(
        n1341) );
  NOR2X1 U72 ( .A(n2891), .B(n2887), .Y(n28) );
  AOI2BB2X1 U73 ( .B0(n2869), .B1(n28), .A0N(n2869), .A1N(n28), .Y(n2894) );
  AO22X1 U74 ( .A0(n29), .A1(n2771), .B0(n2787), .B1(next_work_cntr[5]), .Y(
        n2858) );
  CLKINVX1 U75 ( .A(n2787), .Y(n29) );
  NAND2X1 U76 ( .A(n2139), .B(n1345), .Y(n30) );
  XNOR2X1 U77 ( .A(n30), .B(n933), .Y(n947) );
  NAND2X1 U78 ( .A(n2133), .B(\intadd_3/A[6] ), .Y(n31) );
  AO22X1 U79 ( .A0(n989), .A1(n31), .B0(n994), .B1(n990), .Y(n1003) );
  NAND2BX1 U80 ( .AN(n1879), .B(write_cntr[14]), .Y(n1889) );
  AOI2BB1X1 U81 ( .A0N(n2916), .A1N(n2914), .B0(n2898), .Y(n2912) );
  OAI2BB1X1 U82 ( .A0N(n2375), .A1N(n2671), .B0(n257), .Y(n2650) );
  AOI2BB1X1 U83 ( .A0N(n2499), .A1N(n162), .B0(n2609), .Y(n2624) );
  CLKINVX1 U84 ( .A(n1356), .Y(n33) );
  AOI32X1 U85 ( .A0(n1355), .A1(n33), .A2(n1354), .B0(n1356), .B1(n1359), .Y(
        n1372) );
  OR2X1 U86 ( .A(\DP_OP_725J1_134_142/n202 ), .B(write_addr[9]), .Y(n34) );
  AOI2BB2X1 U87 ( .B0(write_addr[10]), .B1(n34), .A0N(write_addr[10]), .A1N(
        n34), .Y(\DP_OP_725J1_134_142/n260 ) );
  AND2X1 U88 ( .A(write_addr[10]), .B(n34), .Y(\DP_OP_725J1_134_142/n200 ) );
  AO21X1 U89 ( .A0(read_cntr[1]), .A1(read_cntr[0]), .B0(n619), .Y(n709) );
  CLKINVX1 U90 ( .A(n1409), .Y(n35) );
  OAI21XL U91 ( .A0(n1410), .A1(n35), .B0(n777), .Y(n36) );
  AOI2BB1X1 U92 ( .A0N(n208), .A1N(n1409), .B0(n36), .Y(n624) );
  OAI2BB1X1 U93 ( .A0N(n403), .A1N(n404), .B0(n405), .Y(n410) );
  NOR2X1 U94 ( .A(n69), .B(N1453), .Y(n37) );
  AOI211X1 U95 ( .A0(n69), .A1(N1453), .B0(n41), .C0(n37), .Y(n502) );
  AOI21X1 U96 ( .A0(n244), .A1(n2953), .B0(n2952), .Y(next_photo[0]) );
  NOR2X1 U97 ( .A(n814), .B(global_cntr[19]), .Y(n38) );
  AOI211X1 U98 ( .A0(n814), .A1(global_cntr[19]), .B0(n816), .C0(n38), .Y(n782) );
  NOR2BX1 U99 ( .AN(n269), .B(n147), .Y(n39) );
  OA21XL U100 ( .A0(n39), .A1(global_cntr[10]), .B0(n271), .Y(n788) );
  OAI2BB2XL U101 ( .B0(n207), .B1(n42), .A0N(n2945), .A1N(n675), .Y(n493) );
  OA22X1 U102 ( .A0(n2682), .A1(n2681), .B0(n2683), .B1(n2680), .Y(n2728) );
  CLKINVX1 U103 ( .A(n1688), .Y(n74) );
  OR3X2 U104 ( .A(n2499), .B(n162), .C(n146), .Y(n2149) );
  CLKINVX1 U105 ( .A(n2091), .Y(n72) );
  OAI21X1 U106 ( .A0(N2284), .A1(n41), .B0(n2285), .Y(n2299) );
  INVX12 U107 ( .A(reset), .Y(n802) );
  INVX6 U108 ( .A(n42), .Y(n40) );
  OAI21X1 U109 ( .A0(n1690), .A1(n1723), .B0(n1689), .Y(n1699) );
  NAND2X2 U110 ( .A(n1293), .B(n1285), .Y(\next_cr_y[0] ) );
  OAI21X1 U111 ( .A0(n2818), .A1(n2817), .B0(n2816), .Y(n2843) );
  OAI31X1 U112 ( .A0(n984), .A1(n1361), .A2(n983), .B0(n982), .Y(n990) );
  OAI21X1 U113 ( .A0(n2470), .A1(n2469), .B0(n2468), .Y(n2473) );
  NOR2X2 U114 ( .A(n2682), .B(n2677), .Y(n2712) );
  OAI21X1 U115 ( .A0(n1267), .A1(n1266), .B0(n1265), .Y(n1273) );
  OAI21X1 U116 ( .A0(n180), .A1(n1771), .B0(n1770), .Y(n1777) );
  AND2X2 U117 ( .A(n1924), .B(n1922), .Y(n1941) );
  NOR2X1 U118 ( .A(n2546), .B(work_cntr[12]), .Y(n2522) );
  OAI22X1 U119 ( .A0(n1075), .A1(n206), .B0(n1074), .B1(n89), .Y(n1381) );
  NOR2X1 U120 ( .A(n1069), .B(cr_read_cntr[4]), .Y(n503) );
  NOR2X1 U121 ( .A(work_cntr[6]), .B(n2591), .Y(n2576) );
  NAND2X4 U122 ( .A(state[0]), .B(en_so), .Y(n2969) );
  AND2X2 U123 ( .A(state[0]), .B(n281), .Y(n780) );
  NAND2X1 U124 ( .A(curr_time[15]), .B(n1017), .Y(n306) );
  NAND2X1 U125 ( .A(state[0]), .B(n827), .Y(n831) );
  BUFX12 U126 ( .A(n802), .Y(n43) );
  OR4XL U127 ( .A(n781), .B(n2932), .C(n2931), .D(n2930), .Y(n2933) );
  AOI221X1 U128 ( .A0(n2883), .A1(n2882), .B0(n2881), .B1(n2880), .C0(n2879), 
        .Y(n2908) );
  OAI31X1 U129 ( .A0(n2862), .A1(n2865), .A2(n2864), .B0(n2861), .Y(n2900) );
  OAI211X1 U130 ( .A0(n2857), .A1(n2856), .B0(n2855), .C0(n2854), .Y(n2903) );
  AND2X2 U131 ( .A(n108), .B(n109), .Y(n107) );
  NAND2X4 U132 ( .A(n717), .B(n103), .Y(\DP_OP_725J1_134_142/I10 ) );
  NOR2X1 U133 ( .A(n718), .B(n766), .Y(n715) );
  CLKBUFX3 U134 ( .A(n760), .Y(n254) );
  OR2X1 U135 ( .A(n105), .B(n106), .Y(so_mux_sel[0]) );
  OAI31X1 U136 ( .A0(n2295), .A1(n2300), .A2(n2294), .B0(n2293), .Y(n2301) );
  OAI211X1 U137 ( .A0(n1656), .A1(n1655), .B0(n1666), .C0(n1654), .Y(n1679) );
  OAI21X1 U138 ( .A0(n2290), .A1(n2283), .B0(n2282), .Y(n2285) );
  OR2X1 U139 ( .A(n2290), .B(n2279), .Y(n2277) );
  OAI31X1 U140 ( .A0(n972), .A1(n971), .A2(n1361), .B0(n970), .Y(n988) );
  OAI31X1 U141 ( .A0(n1624), .A1(n1614), .A2(n1622), .B0(n1644), .Y(n1643) );
  OAI31X1 U142 ( .A0(n2263), .A1(n2250), .A2(n2257), .B0(n2249), .Y(n2253) );
  OAI21XL U143 ( .A0(n2453), .A1(n2460), .B0(n2454), .Y(n2464) );
  OAI31X1 U144 ( .A0(n942), .A1(n941), .A2(n940), .B0(n939), .Y(n955) );
  OAI31X1 U145 ( .A0(n1144), .A1(n1146), .A2(n1149), .B0(n1143), .Y(n1150) );
  OAI31X1 U146 ( .A0(n1574), .A1(n1565), .A2(n1564), .B0(n61), .Y(n1571) );
  OAI31X1 U147 ( .A0(n130), .A1(n1338), .A2(n1341), .B0(n1337), .Y(n1343) );
  OAI21XL U148 ( .A0(n2433), .A1(n2440), .B0(n2434), .Y(n2444) );
  OA21XL U149 ( .A0(n1834), .A1(n1838), .B0(n1833), .Y(n1840) );
  OA21XL U150 ( .A0(n2424), .A1(n2428), .B0(n2423), .Y(n2431) );
  NOR2X1 U151 ( .A(n1540), .B(n1541), .Y(n1546) );
  OAI31X1 U152 ( .A0(n2081), .A1(n2080), .A2(n2079), .B0(n2078), .Y(n2082) );
  OAI31X1 U153 ( .A0(n904), .A1(n255), .A2(n903), .B0(n902), .Y(n908) );
  OA21XL U154 ( .A0(n1818), .A1(n1822), .B0(n1817), .Y(n1824) );
  OAI31X1 U155 ( .A0(n1813), .A1(work_cntr[6]), .A2(n1812), .B0(n1811), .Y(
        n1820) );
  OAI31X1 U156 ( .A0(n2675), .A1(next_work_cntr[15]), .A2(n2674), .B0(n2673), 
        .Y(n2698) );
  AND3X2 U157 ( .A(n476), .B(n475), .C(n474), .Y(\DP_OP_280J1_126_7605/I3 ) );
  OAI31X1 U158 ( .A0(n889), .A1(n1322), .A2(n888), .B0(n887), .Y(n892) );
  OA21XL U159 ( .A0(n2161), .A1(n2162), .B0(n2176), .Y(n2184) );
  OA21XL U160 ( .A0(n2386), .A1(n2390), .B0(n2385), .Y(n2393) );
  OAI211X1 U161 ( .A0(n2160), .A1(n2163), .B0(n2162), .C0(n2168), .Y(n2176) );
  AOI211X1 U162 ( .A0(n2051), .A1(n2055), .B0(n2050), .C0(n2056), .Y(n2053) );
  OA21XL U163 ( .A0(n1797), .A1(n1796), .B0(n1795), .Y(n1804) );
  OAI31X1 U164 ( .A0(n67), .A1(n1512), .A2(n1511), .B0(n1510), .Y(n1538) );
  AOI31X1 U165 ( .A0(n1943), .A1(n1945), .A2(n1932), .B0(n1948), .Y(n2130) );
  OA21XL U166 ( .A0(n2366), .A1(n2370), .B0(n2365), .Y(n2374) );
  OA22X2 U167 ( .A0(n864), .A1(n2144), .B0(n848), .B1(n847), .Y(n869) );
  OR2X2 U168 ( .A(n132), .B(n133), .Y(n131) );
  CLKAND2X3 U169 ( .A(n257), .B(n2932), .Y(n776) );
  OA21XL U170 ( .A0(n129), .A1(n1252), .B0(n1244), .Y(n1245) );
  OA21XL U171 ( .A0(n1766), .A1(n1770), .B0(n1765), .Y(n1772) );
  OAI31X1 U172 ( .A0(n1761), .A1(work_cntr[12]), .A2(n1760), .B0(n1759), .Y(
        n1768) );
  OAI2BB1X1 U173 ( .A0N(state[0]), .A1N(n837), .B0(n278), .Y(n279) );
  OR2XL U174 ( .A(n1715), .B(n1383), .Y(n1384) );
  OAI222X1 U175 ( .A0(n833), .A1(n2949), .B0(n756), .B1(n830), .C0(n1721), 
        .C1(n2121), .Y(n835) );
  AOI211X1 U176 ( .A0(n148), .A1(n817), .B0(n276), .C0(n816), .Y(n784) );
  OAI31X1 U177 ( .A0(n1745), .A1(n256), .A2(n1744), .B0(n1743), .Y(n1752) );
  OR2XL U178 ( .A(n1388), .B(n1718), .Y(n1389) );
  INVX2 U179 ( .A(n1957), .Y(expand_sel[0]) );
  INVX3 U180 ( .A(n670), .Y(n713) );
  OR2X1 U181 ( .A(n111), .B(n112), .Y(n110) );
  OAI2BB2X2 U182 ( .B0(n129), .B1(n1226), .A0N(n129), .A1N(n1226), .Y(n1246)
         );
  CLKBUFX3 U183 ( .A(n2978), .Y(en_fb_addr) );
  AND2XL U184 ( .A(n286), .B(n294), .Y(n382) );
  OR4XL U185 ( .A(global_cntr[0]), .B(global_cntr[1]), .C(n1954), .D(N2902), 
        .Y(n2979) );
  NOR3X1 U186 ( .A(global_cntr[1]), .B(n183), .C(n1954), .Y(N2880) );
  NOR3X1 U187 ( .A(n1953), .B(n1952), .C(N2902), .Y(n2978) );
  NAND2X1 U188 ( .A(n1873), .B(n150), .Y(n1952) );
  NOR4X1 U189 ( .A(global_cntr[16]), .B(global_cntr[17]), .C(n1872), .D(n1871), 
        .Y(n1873) );
  CLKBUFX3 U190 ( .A(write_addr[13]), .Y(n89) );
  CLKBUFX3 U191 ( .A(write_addr[12]), .Y(n102) );
  BUFX2 U192 ( .A(write_addr[14]), .Y(n88) );
  OAI21X2 U193 ( .A0(work_cntr[18]), .A1(work_cntr[17]), .B0(work_cntr[19]), 
        .Y(n2332) );
  OAI31X1 U194 ( .A0(n2900), .A1(n2889), .A2(n2888), .B0(n2887), .Y(n2890) );
  NAND2X1 U195 ( .A(n2865), .B(n2864), .Y(n2887) );
  CLKINVX1 U196 ( .A(n2464), .Y(n44) );
  CLKINVX1 U197 ( .A(n2444), .Y(n45) );
  NAND2X1 U198 ( .A(n2747), .B(n2746), .Y(n2776) );
  CLKINVX1 U199 ( .A(n382), .Y(n46) );
  NAND2X1 U200 ( .A(n257), .B(n162), .Y(n2284) );
  NOR2BX1 U201 ( .AN(n1933), .B(n1935), .Y(n1936) );
  NAND2X1 U202 ( .A(n806), .B(n198), .Y(n1933) );
  CLKINVX1 U203 ( .A(n1923), .Y(n1935) );
  NAND2X1 U204 ( .A(n310), .B(n319), .Y(n402) );
  BUFX4 U205 ( .A(n613), .Y(n253) );
  NOR2X1 U206 ( .A(n1531), .B(n1530), .Y(n1554) );
  NOR2X1 U207 ( .A(n321), .B(n320), .Y(n368) );
  NOR2X1 U208 ( .A(n318), .B(n317), .Y(n321) );
  NOR2X1 U209 ( .A(n1109), .B(n1304), .Y(n1108) );
  INVXL U210 ( .A(n1384), .Y(n47) );
  OAI2BB2X1 U211 ( .B0(n1986), .B1(n1985), .A0N(n1986), .A1N(n1985), .Y(n1988)
         );
  NOR2X1 U212 ( .A(n2679), .B(next_work_cntr[11]), .Y(n2710) );
  NOR2BX1 U213 ( .AN(n1054), .B(n1301), .Y(n1055) );
  OAI32X1 U214 ( .A0(n2969), .A1(n2325), .A2(n2897), .B0(si_sel), .B1(n2324), 
        .Y(n2927) );
  NAND2X1 U215 ( .A(n2600), .B(n1518), .Y(n1548) );
  NAND2BX1 U216 ( .AN(n1537), .B(n1539), .Y(n1518) );
  NOR2X1 U217 ( .A(n199), .B(n1623), .Y(n1658) );
  CLKINVX1 U218 ( .A(n1201), .Y(n1218) );
  NOR2BX1 U219 ( .AN(\intadd_3/A[0] ), .B(n1301), .Y(n1307) );
  OAI21X1 U220 ( .A0(n193), .A1(n1799), .B0(n1796), .Y(n1793) );
  OAI21X1 U221 ( .A0(n150), .A1(n1874), .B0(n2321), .Y(n834) );
  OAI211X1 U222 ( .A0(n479), .A1(n241), .B0(cr_read_cntr[3]), .C0(n477), .Y(
        n505) );
  NOR2X1 U223 ( .A(n137), .B(n173), .Y(n1416) );
  NOR2BX1 U224 ( .AN(n2509), .B(work_cntr[19]), .Y(n2513) );
  NOR2BX1 U225 ( .AN(next_cr_x[6]), .B(n1304), .Y(n1309) );
  INVX3 U226 ( .A(n1305), .Y(n1304) );
  OAI21X1 U227 ( .A0(n2341), .A1(n2340), .B0(n2339), .Y(n2349) );
  INVXL U228 ( .A(n2393), .Y(n49) );
  OAI21X1 U229 ( .A0(n1750), .A1(n1754), .B0(n1749), .Y(n1757) );
  OAI21X1 U230 ( .A0(n2347), .A1(n2351), .B0(n2346), .Y(n2355) );
  INVXL U231 ( .A(n2374), .Y(n50) );
  OAI21X1 U232 ( .A0(n2955), .A1(n1865), .B0(n2963), .Y(n1864) );
  OAI21X1 U233 ( .A0(n1734), .A1(n1733), .B0(n1732), .Y(n1740) );
  INVXL U234 ( .A(n1824), .Y(n51) );
  INVXL U235 ( .A(n1840), .Y(n52) );
  INVXL U236 ( .A(n2431), .Y(n53) );
  INVXL U237 ( .A(n1804), .Y(n54) );
  OAI21X1 U238 ( .A0(n1802), .A1(n1806), .B0(n1801), .Y(n1808) );
  OAI21X1 U239 ( .A0(n2404), .A1(n2408), .B0(n2403), .Y(n2411) );
  AOI32X1 U240 ( .A0(n1731), .A1(n1730), .A2(n181), .B0(n1738), .B1(n1730), 
        .Y(n1736) );
  NOR2X1 U241 ( .A(n1729), .B(n1728), .Y(n1738) );
  CLKINVX1 U242 ( .A(n1544), .Y(n1552) );
  NAND2X1 U243 ( .A(n862), .B(n861), .Y(n1058) );
  NAND2X1 U244 ( .A(n862), .B(n860), .Y(n861) );
  OAI21X1 U245 ( .A0(n928), .A1(n927), .B0(n926), .Y(n937) );
  OAI2BB1X1 U246 ( .A0N(n1961), .A1N(work_cntr[17]), .B0(n1963), .Y(n1982) );
  NAND3X1 U247 ( .A(n2014), .B(n1960), .C(n182), .Y(n1963) );
  OAI21X1 U248 ( .A0(n1132), .A1(n1131), .B0(n1130), .Y(n1152) );
  OAI21X1 U249 ( .A0(n2794), .A1(n2793), .B0(n2792), .Y(n2815) );
  OAI2BB2X1 U250 ( .B0(n1343), .B1(n1342), .A0N(n1343), .A1N(n1345), .Y(n1353)
         );
  AND2X2 U251 ( .A(n1346), .B(n1345), .Y(n1342) );
  INVX3 U252 ( .A(n940), .Y(n1345) );
  INVXL U253 ( .A(n1772), .Y(n55) );
  NOR2X2 U254 ( .A(n165), .B(n146), .Y(n2120) );
  OAI21X1 U255 ( .A0(work_cntr[4]), .A1(n41), .B0(n2278), .Y(n2286) );
  NOR2X1 U256 ( .A(n2820), .B(n2819), .Y(n2849) );
  OAI2BB2X1 U257 ( .B0(n2144), .B1(n1877), .A0N(n2144), .A1N(n1877), .Y(n1882)
         );
  AOI2BB2X2 U258 ( .B0(n2142), .B1(n1053), .A0N(n2142), .A1N(n1053), .Y(n1096)
         );
  OAI21X1 U259 ( .A0(n2619), .A1(n2618), .B0(n2617), .Y(n2623) );
  AOI2BB2X2 U260 ( .B0(n2533), .B1(n2532), .A0N(n2533), .A1N(n2531), .Y(n2544)
         );
  OAI22X1 U261 ( .A0(write_addr[9]), .A1(n1367), .B0(n233), .B1(n1366), .Y(
        n1370) );
  INVXL U262 ( .A(N633), .Y(n56) );
  INVXL U263 ( .A(n56), .Y(n57) );
  OAI21X1 U264 ( .A0(n973), .A1(n907), .B0(n864), .Y(n906) );
  INVX3 U265 ( .A(n131), .Y(n973) );
  OAI22X1 U266 ( .A0(n885), .A1(n884), .B0(n883), .B1(n882), .Y(n896) );
  OAI22X1 U267 ( .A0(n2502), .A1(n2521), .B0(n256), .B1(n2503), .Y(n2538) );
  NOR3X1 U268 ( .A(n2615), .B(n2614), .C(n2613), .Y(n2621) );
  INVXL U269 ( .A(n2466), .Y(n58) );
  INVXL U270 ( .A(n58), .Y(n59) );
  OAI31X1 U271 ( .A0(n900), .A1(n899), .A2(n255), .B0(n898), .Y(n914) );
  XOR2X1 U272 ( .A(\DP_OP_725J1_134_142/n146 ), .B(\DP_OP_725J1_134_142/n145 ), 
        .Y(N1686) );
  AND2X2 U273 ( .A(n2761), .B(n2762), .Y(n2736) );
  INVXL U274 ( .A(n1572), .Y(n60) );
  INVXL U275 ( .A(n60), .Y(n61) );
  OAI31X1 U276 ( .A0(n2045), .A1(n2044), .A2(n2043), .B0(n2042), .Y(n2046) );
  AOI2BB2X2 U277 ( .B0(work_cntr[13]), .B1(n1202), .A0N(work_cntr[13]), .A1N(
        n1202), .Y(n1206) );
  NOR2X1 U278 ( .A(n233), .B(n1369), .Y(n1368) );
  OAI21X2 U279 ( .A0(n1683), .A1(write_addr[8]), .B0(n1366), .Y(n1369) );
  NOR2BX1 U280 ( .AN(n1453), .B(n161), .Y(n1447) );
  OAI31X1 U281 ( .A0(n1475), .A1(n1474), .A2(n1486), .B0(n1473), .Y(n1523) );
  NOR2X1 U282 ( .A(work_cntr[13]), .B(n1501), .Y(n1475) );
  NOR2BX1 U283 ( .AN(n2052), .B(n2051), .Y(n2062) );
  NAND2X2 U284 ( .A(im_wen_n), .B(n257), .Y(n2945) );
  CLKINVX1 U285 ( .A(n2152), .Y(n2217) );
  OAI22X2 U286 ( .A0(n2684), .A1(n2217), .B0(next_work_cntr[11]), .B1(n2152), 
        .Y(n2216) );
  NOR2X1 U287 ( .A(n2218), .B(next_work_cntr[10]), .Y(n2152) );
  NOR2X1 U288 ( .A(next_work_cntr[6]), .B(n2252), .Y(n2150) );
  NAND2X1 U289 ( .A(curr_time[7]), .B(n1024), .Y(n319) );
  NOR2X1 U290 ( .A(curr_time[10]), .B(n392), .Y(n441) );
  XOR2X1 U291 ( .A(n402), .B(curr_time[4]), .Y(n1026) );
  AND2X2 U292 ( .A(n1630), .B(n1625), .Y(n1637) );
  NAND2X1 U293 ( .A(n199), .B(n1623), .Y(n1657) );
  CLKINVX1 U294 ( .A(n446), .Y(n434) );
  AND3X2 U295 ( .A(n395), .B(n394), .C(n393), .Y(n446) );
  NOR2X1 U296 ( .A(n2077), .B(n2084), .Y(n2079) );
  NAND2X1 U297 ( .A(n2076), .B(n164), .Y(n2084) );
  OAI31X1 U298 ( .A0(n2438), .A1(n2437), .A2(n2436), .B0(n2435), .Y(n2446) );
  NAND2X1 U299 ( .A(n2427), .B(n2429), .Y(n2438) );
  OAI31X1 U300 ( .A0(n1829), .A1(work_cntr[4]), .A2(n1828), .B0(n1827), .Y(
        n1836) );
  NAND2X1 U301 ( .A(n1821), .B(n1823), .Y(n1829) );
  OAI31X1 U302 ( .A0(n2418), .A1(n2417), .A2(n2416), .B0(n2415), .Y(n2426) );
  NAND2X1 U303 ( .A(n2407), .B(n2409), .Y(n2418) );
  OAI31X1 U304 ( .A0(n2398), .A1(n2649), .A2(n2397), .B0(n2396), .Y(n2406) );
  NAND2X1 U305 ( .A(n2389), .B(n2391), .Y(n2398) );
  OAI31X1 U306 ( .A0(n2380), .A1(n2379), .A2(n2378), .B0(n2377), .Y(n2388) );
  NAND2X1 U307 ( .A(n2369), .B(n2371), .Y(n2380) );
  NAND2X1 U308 ( .A(n1753), .B(n1755), .Y(n1761) );
  OAI31X1 U309 ( .A0(n2361), .A1(n2360), .A2(n2359), .B0(n2358), .Y(n2368) );
  NAND2X1 U310 ( .A(n2350), .B(n2352), .Y(n2361) );
  NAND2X1 U311 ( .A(n1805), .B(n1807), .Y(n1813) );
  NAND2X1 U312 ( .A(n881), .B(n1052), .Y(n1054) );
  NOR2X1 U313 ( .A(n2135), .B(n1093), .Y(n1052) );
  NAND2X1 U314 ( .A(n1650), .B(n1661), .Y(n1665) );
  OAI211X1 U315 ( .A0(n1663), .A1(n1662), .B0(n1661), .C0(n1664), .Y(n1678) );
  CLKINVX1 U316 ( .A(n1624), .Y(n1661) );
  NAND2X1 U317 ( .A(n796), .B(global_cntr[3]), .Y(n263) );
  OA21X2 U318 ( .A0(n1289), .A1(\intadd_3/A[0] ), .B0(n1288), .Y(n1411) );
  OAI31X1 U319 ( .A0(n175), .A1(n867), .A2(n1321), .B0(n868), .Y(n886) );
  CLKINVX1 U320 ( .A(n870), .Y(n1321) );
  CLKINVX1 U321 ( .A(n995), .Y(n1007) );
  AND3X2 U322 ( .A(n69), .B(N1453), .C(N1454), .Y(n359) );
  NOR2X2 U323 ( .A(n2059), .B(n2058), .Y(n2075) );
  CLKINVX1 U324 ( .A(n1849), .Y(n1853) );
  NAND2X1 U325 ( .A(n1843), .B(n1842), .Y(n1849) );
  CLKINVX1 U326 ( .A(n2375), .Y(n2379) );
  NOR2X1 U327 ( .A(n197), .B(n1543), .Y(n1567) );
  NOR2BX1 U328 ( .AN(n1566), .B(n1567), .Y(n1597) );
  NAND2X1 U329 ( .A(n197), .B(n1543), .Y(n1566) );
  NOR2X1 U330 ( .A(n2190), .B(n2196), .Y(n2200) );
  NAND2X1 U331 ( .A(n2190), .B(n2189), .Y(n2209) );
  NAND2X1 U332 ( .A(n2180), .B(n2179), .Y(n2189) );
  CLKINVX1 U333 ( .A(n2587), .Y(n2594) );
  NAND2X1 U334 ( .A(n1450), .B(n182), .Y(n1724) );
  CLKINVX1 U335 ( .A(n2356), .Y(n2360) );
  CLKINVX1 U336 ( .A(n2867), .Y(n2865) );
  AOI2BB2X2 U337 ( .B0(next_work_cntr[6]), .B1(n2252), .A0N(next_work_cntr[6]), 
        .A1N(n2252), .Y(n2265) );
  OAI31X4 U338 ( .A0(n68), .A1(n164), .A2(n41), .B0(n2771), .Y(n2252) );
  NOR2X1 U339 ( .A(n1348), .B(n1135), .Y(n949) );
  NAND2X1 U340 ( .A(n872), .B(n882), .Y(n888) );
  NAND2X1 U341 ( .A(n885), .B(n2142), .Y(n882) );
  NAND2X1 U342 ( .A(n424), .B(n416), .Y(n425) );
  AOI31X1 U343 ( .A0(n1013), .A1(curr_time[18]), .A2(n410), .B0(n406), .Y(n424) );
  NOR2X1 U344 ( .A(n1458), .B(n1470), .Y(n1461) );
  NAND2X1 U345 ( .A(n187), .B(n1457), .Y(n1470) );
  NOR2X1 U346 ( .A(n2109), .B(n2969), .Y(expand_sel[3]) );
  AND2X2 U347 ( .A(n2082), .B(N2284), .Y(n2090) );
  NAND2X1 U348 ( .A(n2731), .B(n2730), .Y(n2724) );
  NAND2X1 U349 ( .A(n1735), .B(n1736), .Y(n1739) );
  NAND2X1 U350 ( .A(N2283), .B(N2282), .Y(n2499) );
  NOR2X1 U351 ( .A(n2027), .B(n2026), .Y(n2033) );
  AOI31X1 U352 ( .A0(n2866), .A1(n2884), .A2(n2886), .B0(n2894), .Y(n2893) );
  NOR2X1 U353 ( .A(n2900), .B(n2911), .Y(n2886) );
  NOR2X1 U354 ( .A(n2764), .B(n2765), .Y(n2755) );
  NAND2X1 U355 ( .A(n2735), .B(n2752), .Y(n2765) );
  NAND2X1 U356 ( .A(n193), .B(n1488), .Y(n1504) );
  NAND2BX1 U357 ( .AN(n1468), .B(n1467), .Y(n1488) );
  NOR2X1 U358 ( .A(n2172), .B(n76), .Y(n2182) );
  NOR2BX1 U359 ( .AN(n1488), .B(n1487), .Y(n1492) );
  NAND2X1 U360 ( .A(n896), .B(n895), .Y(n903) );
  NAND2X1 U361 ( .A(n894), .B(n2141), .Y(n895) );
  CLKINVX1 U362 ( .A(n2795), .Y(next_work_cntr[4]) );
  NAND2X1 U363 ( .A(n257), .B(n2457), .Y(n2795) );
  NAND2X1 U364 ( .A(n1723), .B(n1722), .Y(n2113) );
  NOR2X1 U365 ( .A(n75), .B(n2966), .Y(n1723) );
  NOR2X1 U366 ( .A(n2934), .B(n240), .Y(n2935) );
  NOR2X1 U367 ( .A(n2939), .B(n242), .Y(n2940) );
  NAND2X1 U368 ( .A(n2132), .B(n999), .Y(n1000) );
  NOR2BX1 U369 ( .AN(\s_1[2] ), .B(curr_time[3]), .Y(n1027) );
  NAND2X1 U370 ( .A(n369), .B(n368), .Y(\s_1[2] ) );
  NOR2BX1 U371 ( .AN(n2898), .B(n2911), .Y(n2877) );
  NOR2X1 U372 ( .A(n1700), .B(n772), .Y(n1711) );
  NAND2X1 U373 ( .A(n1706), .B(n1721), .Y(n1700) );
  NOR2X1 U374 ( .A(n2484), .B(n2483), .Y(n2487) );
  OAI21X1 U375 ( .A0(n1121), .A1(n1134), .B0(n1120), .Y(n1122) );
  NAND2X1 U376 ( .A(n1135), .B(\intadd_3/A[0] ), .Y(n1134) );
  NOR2X1 U377 ( .A(n1998), .B(n1997), .Y(n2004) );
  OAI21X1 U378 ( .A0(n2487), .A1(n2485), .B0(n2486), .Y(n2490) );
  NOR2BX1 U379 ( .AN(n2481), .B(n2475), .Y(n2485) );
  NOR2X1 U380 ( .A(n2216), .B(n2215), .Y(n2214) );
  NOR2X1 U381 ( .A(N2282), .B(n41), .Y(n2305) );
  NAND2X1 U382 ( .A(n2771), .B(n2787), .Y(n2829) );
  NAND2X1 U383 ( .A(n1000), .B(n1003), .Y(n1006) );
  NAND2X1 U384 ( .A(n257), .B(n2442), .Y(n2771) );
  NOR2X1 U385 ( .A(n2225), .B(n2224), .Y(n2208) );
  NAND2X1 U386 ( .A(n2027), .B(n2026), .Y(n2037) );
  NOR2X1 U387 ( .A(n1865), .B(n1963), .Y(n1166) );
  NOR2X2 U388 ( .A(next_work_cntr[2]), .B(n2863), .Y(n2876) );
  OAI2BB2X2 U389 ( .B0(next_work_cntr[2]), .B1(n2863), .A0N(next_work_cntr[2]), 
        .A1N(n2863), .Y(n2911) );
  AND2X2 U390 ( .A(n2847), .B(n2873), .Y(n2863) );
  NOR2BX1 U391 ( .AN(n1713), .B(n1369), .Y(n1362) );
  OAI21X1 U392 ( .A0(work_cntr[19]), .A1(n1168), .B0(n1167), .Y(n1172) );
  AOI211X1 U393 ( .A0(n1962), .A1(n1254), .B0(n1168), .C0(n152), .Y(n1169) );
  NOR2X1 U394 ( .A(n1166), .B(n161), .Y(n1168) );
  OAI31X1 U395 ( .A0(n2276), .A1(n2275), .A2(n2274), .B0(n2273), .Y(n2278) );
  NOR2X1 U396 ( .A(n2280), .B(n2279), .Y(n2274) );
  AOI21X1 U397 ( .A0(n2671), .A1(n2678), .B0(n2670), .Y(n2677) );
  NAND2X1 U398 ( .A(n257), .B(n2379), .Y(n2670) );
  NAND2X1 U399 ( .A(global_cntr[7]), .B(n266), .Y(n267) );
  NAND2X1 U400 ( .A(global_cntr[16]), .B(n273), .Y(n817) );
  NAND2BX1 U401 ( .AN(n1647), .B(n1668), .Y(n1646) );
  NOR2X1 U402 ( .A(n2169), .B(n2170), .Y(n2181) );
  NOR2X1 U403 ( .A(n296), .B(n295), .Y(n404) );
  NAND2X1 U404 ( .A(n2932), .B(n2322), .Y(n2950) );
  CLKINVX1 U405 ( .A(n1456), .Y(n1494) );
  NOR2BX1 U406 ( .AN(n2196), .B(n2195), .Y(n2204) );
  NOR2X1 U407 ( .A(n2179), .B(n2180), .Y(n2195) );
  NOR2X1 U408 ( .A(n1335), .B(n1057), .Y(n912) );
  OAI31X1 U409 ( .A0(n1279), .A1(n1280), .A2(n2486), .B0(n1277), .Y(n2959) );
  NOR2X1 U410 ( .A(n2476), .B(n1276), .Y(n1280) );
  NOR2X1 U411 ( .A(n1993), .B(n2002), .Y(n2007) );
  AOI32X1 U412 ( .A0(n839), .A1(n838), .A2(n854), .B0(n189), .B1(n838), .Y(
        n2930) );
  NOR2X1 U413 ( .A(write_cntr[9]), .B(write_cntr[10]), .Y(n839) );
  NOR2X1 U414 ( .A(n2102), .B(n2101), .Y(n2106) );
  NAND2X1 U415 ( .A(global_cntr[12]), .B(n270), .Y(n259) );
  AOI31X1 U416 ( .A0(n911), .A1(n910), .A2(n1334), .B0(n909), .Y(n928) );
  NAND2X1 U417 ( .A(n2135), .B(n913), .Y(n911) );
  NOR2X1 U418 ( .A(n2836), .B(n2835), .Y(n2814) );
  NOR2BX1 U419 ( .AN(n1542), .B(n1536), .Y(n1540) );
  NOR2BX1 U420 ( .AN(n1704), .B(n1721), .Y(n1695) );
  NOR2X1 U421 ( .A(n1103), .B(n2140), .Y(n1091) );
  NOR2X1 U422 ( .A(n1866), .B(n146), .Y(n2960) );
  NAND2X1 U423 ( .A(n165), .B(n1646), .Y(n1673) );
  OAI21X1 U424 ( .A0(n1658), .A1(n1673), .B0(n1657), .Y(n1659) );
  OAI21X1 U425 ( .A0(n2236), .A1(n2220), .B0(n2219), .Y(n2231) );
  NAND2BX1 U426 ( .AN(n2222), .B(n2224), .Y(n2220) );
  OAI2BB2X1 U427 ( .B0(n2554), .B1(n2553), .A0N(n2554), .A1N(n2556), .Y(n2558)
         );
  NOR2BX1 U428 ( .AN(n1495), .B(n1517), .Y(n1515) );
  OAI2BB2X1 U429 ( .B0(n1494), .B1(n1493), .A0N(n1494), .A1N(n1493), .Y(n1517)
         );
  NOR2BX1 U430 ( .AN(n1623), .B(n1622), .Y(n1653) );
  NAND2X1 U431 ( .A(n184), .B(n2522), .Y(n2521) );
  NOR2BX1 U432 ( .AN(n2530), .B(n2520), .Y(n2535) );
  AOI21X2 U433 ( .A0(n2600), .A1(n1045), .B0(n1044), .Y(n2437) );
  NAND2BX1 U434 ( .AN(n994), .B(n993), .Y(n987) );
  NOR2BX1 U435 ( .AN(n1581), .B(n1580), .Y(n1632) );
  NOR2X1 U436 ( .A(n206), .B(n1380), .Y(n1387) );
  AOI21X2 U437 ( .A0(n188), .A1(n1035), .B0(n1034), .Y(n2660) );
  AOI21X1 U438 ( .A0(n1539), .A1(n1538), .B0(n1537), .Y(n1541) );
  AOI31X1 U439 ( .A0(n1551), .A1(n1514), .A2(n81), .B0(n1538), .Y(n1537) );
  NOR2X1 U440 ( .A(n1651), .B(n1673), .Y(n1663) );
  NOR2X1 U441 ( .A(n1304), .B(n1296), .Y(\intadd_3/B[0] ) );
  OAI21X1 U442 ( .A0(n1295), .A1(n1294), .B0(n1293), .Y(n1296) );
  OAI21X1 U443 ( .A0(n2328), .A1(n2329), .B0(n2327), .Y(n2335) );
  AOI221X1 U444 ( .A0(n948), .A1(n947), .B0(n946), .B1(n947), .C0(n954), .Y(
        n963) );
  NOR2X1 U445 ( .A(n1348), .B(n945), .Y(n954) );
  OAI2BB2X1 U446 ( .B0(n2284), .B1(n2285), .A0N(n2284), .A1N(n2285), .Y(n2294)
         );
  OAI21X1 U447 ( .A0(n165), .A1(n1852), .B0(n1857), .Y(n1858) );
  OAI21X1 U448 ( .A0(n2745), .A1(n2744), .B0(n2743), .Y(n2767) );
  NAND2X1 U449 ( .A(n1643), .B(n1642), .Y(n1623) );
  OAI21X1 U450 ( .A0(n1618), .A1(n1617), .B0(n1616), .Y(n1642) );
  OAI21X1 U451 ( .A0(n45), .A1(n2448), .B0(n2443), .Y(n2452) );
  OAI21X1 U452 ( .A0(n2851), .A1(n2876), .B0(n2850), .Y(n2852) );
  AND2X2 U453 ( .A(n2819), .B(n2820), .Y(n2851) );
  NAND2X1 U454 ( .A(n1479), .B(n180), .Y(n1458) );
  OAI21X1 U455 ( .A0(n1853), .A1(n1851), .B0(n165), .Y(n1857) );
  CLKINVX1 U456 ( .A(n2555), .Y(n2567) );
  OAI21X1 U457 ( .A0(n2559), .A1(n180), .B0(n2546), .Y(n2555) );
  AOI211X4 U458 ( .A0(n140), .A1(n274), .B0(n275), .C0(n816), .Y(n785) );
  CLKINVX1 U459 ( .A(n2537), .Y(n2550) );
  OAI21X1 U460 ( .A0(n2522), .A1(n184), .B0(n2521), .Y(n2537) );
  CLKINVX1 U461 ( .A(n1251), .Y(n1259) );
  OAI21X1 U462 ( .A0(n1243), .A1(n197), .B0(n1242), .Y(n1251) );
  AOI22X1 U463 ( .A0(n2585), .A1(n2584), .B0(n2583), .B1(n2582), .Y(n2589) );
  OAI21X1 U464 ( .A0(n2580), .A1(n2579), .B0(n2578), .Y(n2585) );
  CLKINVX1 U465 ( .A(n2610), .Y(n2615) );
  AOI22X1 U466 ( .A0(n2612), .A1(n2611), .B0(n2614), .B1(n2610), .Y(n2620) );
  OAI21X1 U467 ( .A0(n2592), .A1(n197), .B0(n2591), .Y(n2610) );
  CLKINVX1 U468 ( .A(n2066), .Y(n2074) );
  OAI21X1 U469 ( .A0(n2057), .A1(n2059), .B0(n2058), .Y(n2066) );
  OAI21X1 U470 ( .A0(n1935), .A1(n1934), .B0(n1933), .Y(n1940) );
  NOR2X1 U471 ( .A(cr_read_cntr[8]), .B(n237), .Y(n1064) );
  NAND2X1 U472 ( .A(global_cntr[14]), .B(n260), .Y(n272) );
  AND2X2 U473 ( .A(global_cntr[1]), .B(global_cntr[0]), .Y(n798) );
  NAND2X1 U474 ( .A(global_cntr[1]), .B(n183), .Y(n1874) );
  NOR2X1 U475 ( .A(n238), .B(n1068), .Y(n1066) );
  OAI21X1 U476 ( .A0(cr_read_cntr[6]), .A1(n1064), .B0(n1063), .Y(n1068) );
  AOI211X1 U477 ( .A0(n238), .A1(n1068), .B0(n1067), .C0(n1066), .Y(n1071) );
  NAND2X1 U478 ( .A(n257), .B(n2437), .Y(n2751) );
  NOR2X1 U479 ( .A(n2472), .B(n2471), .Y(n2475) );
  OAI21X1 U480 ( .A0(n44), .A1(n2468), .B0(n2463), .Y(n2472) );
  OAI2BB2X1 U481 ( .B0(n1533), .B1(n1476), .A0N(n1533), .A1N(n1476), .Y(n1532)
         );
  NOR2X2 U482 ( .A(n2754), .B(n2775), .Y(n2807) );
  NOR2X1 U483 ( .A(n2751), .B(n2750), .Y(n2775) );
  NOR2X1 U484 ( .A(n1773), .B(n55), .Y(n1775) );
  OAI22X1 U485 ( .A0(n1375), .A1(n1374), .B0(n1373), .B1(n1372), .Y(
        \intadd_3/A[8] ) );
  NAND2X1 U486 ( .A(n1375), .B(n1374), .Y(n1373) );
  OAI211X1 U487 ( .A0(n1360), .A1(n1359), .B0(n1358), .C0(n1357), .Y(n1374) );
  OAI211X1 U488 ( .A0(n2638), .A1(n2639), .B0(n2637), .C0(n2636), .Y(n2643) );
  NAND2X1 U489 ( .A(n2970), .B(n2969), .Y(so_mux_sel[1]) );
  OAI21X1 U490 ( .A0(n1416), .A1(N744), .B0(n1424), .Y(n1422) );
  AOI2BB2X2 U491 ( .B0(n1093), .B1(n1092), .A0N(n1093), .A1N(n1092), .Y(n1110)
         );
  OAI21X1 U492 ( .A0(n2135), .A1(n1301), .B0(n1106), .Y(n1092) );
  CLKINVX1 U493 ( .A(n2499), .Y(n2629) );
  NOR2X1 U494 ( .A(n1080), .B(n136), .Y(n1079) );
  AOI2BB2X2 U495 ( .B0(n2588), .B1(n2587), .A0N(n2588), .A1N(n2586), .Y(n2596)
         );
  OAI21X1 U496 ( .A0(n2574), .A1(n2582), .B0(n2590), .Y(n2588) );
  OAI211X1 U497 ( .A0(n772), .A1(write_addr[8]), .B0(n1703), .C0(n1702), .Y(
        n1707) );
  OAI21X1 U498 ( .A0(n2479), .A1(n2480), .B0(n2478), .Y(n2484) );
  OAI21X1 U499 ( .A0(n2475), .A1(n2474), .B0(n2482), .Y(n2480) );
  OAI21X1 U500 ( .A0(n1213), .A1(n1212), .B0(n1225), .Y(n1224) );
  OAI21X1 U501 ( .A0(n1781), .A1(n1780), .B0(n1779), .Y(n1787) );
  OAI21X1 U502 ( .A0(n1775), .A1(n1774), .B0(n160), .Y(n1780) );
  AOI21X1 U503 ( .A0(n1582), .A1(n1583), .B0(n1584), .Y(n1609) );
  OAI211X1 U504 ( .A0(n1579), .A1(n1578), .B0(n1577), .C0(n1576), .Y(n1583) );
  OAI21X1 U505 ( .A0(n1549), .A1(n1566), .B0(n1548), .Y(n1550) );
  NOR2X1 U506 ( .A(n2600), .B(n1518), .Y(n1549) );
  OAI31X1 U507 ( .A0(n1142), .A1(n2137), .A2(n1141), .B0(n1140), .Y(n1147) );
  OAI21X1 U508 ( .A0(\intadd_3/A[0] ), .A1(n1135), .B0(n1134), .Y(n1142) );
  OAI22X1 U509 ( .A0(n2572), .A1(n2580), .B0(n2571), .B1(n2570), .Y(n2581) );
  NAND2X1 U510 ( .A(n264), .B(global_cntr[5]), .Y(n818) );
  OAI22X1 U511 ( .A0(n2781), .A1(n2780), .B0(n2779), .B1(n2791), .Y(n2817) );
  OAI31X1 U512 ( .A0(n2003), .A1(n2002), .A2(n2001), .B0(n2000), .Y(n2008) );
  AOI21X1 U513 ( .A0(n2000), .A1(n1994), .B0(n1993), .Y(n1998) );
  OAI221X1 U514 ( .A0(n1997), .A1(n1990), .B0(n2006), .B1(n1990), .C0(n2003), 
        .Y(n2000) );
  OAI22X1 U515 ( .A0(n1137), .A1(n1136), .B0(n1135), .B1(\intadd_3/A[0] ), .Y(
        n1138) );
  NOR3BX1 U516 ( .AN(n1139), .B(n1142), .C(n2134), .Y(n1144) );
  NAND3X1 U517 ( .A(n1139), .B(n1123), .C(n1135), .Y(n1124) );
  OAI22X2 U518 ( .A0(n1119), .A1(n1304), .B0(n2139), .B1(n1305), .Y(n1139) );
  NAND3X1 U519 ( .A(write_cntr[1]), .B(write_cntr[0]), .C(write_cntr[2]), .Y(
        n931) );
  NOR2X1 U520 ( .A(n2178), .B(n2181), .Y(n2172) );
  NOR3X1 U521 ( .A(n2169), .B(n76), .C(n2171), .Y(n2178) );
  OAI22X1 U522 ( .A0(n1050), .A1(n1049), .B0(n1058), .B1(n1048), .Y(n1099) );
  NOR2X1 U523 ( .A(n2227), .B(n2214), .Y(n2236) );
  NOR2X1 U524 ( .A(n2227), .B(n2226), .Y(n2229) );
  NOR3X1 U525 ( .A(n2216), .B(n2225), .C(n2220), .Y(n2227) );
  NOR3X1 U526 ( .A(write_cntr[14]), .B(write_cntr[12]), .C(write_cntr[13]), 
        .Y(n838) );
  AOI31X4 U527 ( .A0(n2056), .A1(n2055), .A2(n2054), .B0(n2053), .Y(n2059) );
  OAI31X1 U528 ( .A0(n880), .A1(n879), .A2(n1322), .B0(n878), .Y(n901) );
  OAI31X1 U529 ( .A0(n917), .A1(n1335), .A2(n916), .B0(n915), .Y(n919) );
  NOR2X1 U530 ( .A(n2088), .B(n2087), .Y(n2104) );
  NOR3X1 U531 ( .A(n162), .B(n2077), .C(n72), .Y(n2088) );
  NOR3BX1 U532 ( .AN(n1246), .B(n1247), .C(n1244), .Y(n1253) );
  AOI21X1 U533 ( .A0(n1257), .A1(n1256), .B0(n1255), .Y(n1261) );
  NOR3X1 U534 ( .A(n1256), .B(n1253), .C(n1257), .Y(n1255) );
  CLKINVX1 U535 ( .A(n2737), .Y(n2758) );
  NOR3X2 U536 ( .A(n785), .B(n784), .C(n824), .Y(n2321) );
  NAND2X1 U537 ( .A(n1150), .B(n1152), .Y(n1299) );
  AOI2BB2X2 U538 ( .B0(n2838), .B1(n2837), .A0N(n2838), .A1N(n2837), .Y(n2869)
         );
  AOI2BB2X2 U539 ( .B0(n2552), .B1(n2551), .A0N(n2552), .A1N(n2550), .Y(n2564)
         );
  OAI21X1 U540 ( .A0(n2565), .A1(n2564), .B0(n2563), .Y(n2569) );
  AOI2BB2X2 U541 ( .B0(n2569), .B1(n2568), .A0N(n2569), .A1N(n2567), .Y(n2579)
         );
  AOI2BB2X2 U542 ( .B0(n1534), .B1(n1533), .A0N(n1534), .A1N(n1532), .Y(n1592)
         );
  NOR2X1 U543 ( .A(n2836), .B(n2825), .Y(n2808) );
  NOR2X1 U544 ( .A(n2825), .B(n2832), .Y(n2810) );
  AOI2BB2X2 U545 ( .B0(n2773), .B1(n2822), .A0N(n2773), .A1N(n2822), .Y(n2825)
         );
  NAND2BX1 U546 ( .AN(n2932), .B(n781), .Y(n2926) );
  NOR2X2 U547 ( .A(next_state[2]), .B(next_state[1]), .Y(n2932) );
  OAI211X1 U548 ( .A0(n87), .A1(n1686), .B0(n1689), .C0(n1681), .Y(n1722) );
  NOR4X1 U549 ( .A(n1680), .B(n1679), .C(n1678), .D(n1677), .Y(n1689) );
  CLKINVX1 U550 ( .A(n2979), .Y(en_photo_num) );
  NOR2X1 U551 ( .A(N2284), .B(n2955), .Y(n2644) );
  OA21XL U552 ( .A0(n208), .A1(n1083), .B0(n1683), .Y(n1087) );
  NAND4X1 U553 ( .A(N2283), .B(N205), .C(n2644), .D(n165), .Y(n2962) );
  AOI21X1 U554 ( .A0(n142), .A1(n267), .B0(n269), .Y(n790) );
  OAI21X1 U555 ( .A0(n936), .A1(n935), .B0(n934), .Y(n943) );
  NOR2X1 U556 ( .A(n941), .B(n942), .Y(n936) );
  AND2X2 U557 ( .A(n2727), .B(n2726), .Y(n2762) );
  NOR2X1 U558 ( .A(n2720), .B(n2724), .Y(n2726) );
  AOI211X1 U559 ( .A0(n2508), .A1(work_cntr[19]), .B0(n2509), .C0(n2507), .Y(
        n2510) );
  NOR2X1 U560 ( .A(n2505), .B(work_cntr[18]), .Y(n2508) );
  NOR2X1 U561 ( .A(n256), .B(n1959), .Y(n1967) );
  OAI21X1 U562 ( .A0(n1967), .A1(n188), .B0(n1966), .Y(n1971) );
  NOR2X1 U563 ( .A(n2857), .B(n2848), .Y(n2870) );
  NOR2BX1 U564 ( .AN(n1988), .B(n1987), .Y(n2002) );
  AOI21X1 U565 ( .A0(n256), .A1(n1959), .B0(n1967), .Y(n1987) );
  NOR3X1 U566 ( .A(n1987), .B(n1989), .C(n1992), .Y(n1993) );
  NAND2BX1 U567 ( .AN(n1988), .B(n1987), .Y(n2006) );
  NOR2X1 U568 ( .A(n2806), .B(n2853), .Y(n2831) );
  NOR2X1 U569 ( .A(n2707), .B(n2704), .Y(n2722) );
  NOR2X1 U570 ( .A(n2830), .B(n2827), .Y(n2826) );
  OAI2BB1X2 U571 ( .A0N(n386), .A1N(n385), .B0(n384), .Y(n440) );
  NAND2X1 U572 ( .A(n384), .B(n386), .Y(m_1[2]) );
  NOR2X1 U573 ( .A(n308), .B(n307), .Y(n386) );
  NAND2X1 U574 ( .A(n1606), .B(n1605), .Y(n1649) );
  NOR2X1 U575 ( .A(n1596), .B(n1626), .Y(n1606) );
  OAI221X1 U576 ( .A0(n1605), .A1(n1606), .B0(n1602), .B1(n1601), .C0(n1600), 
        .Y(n1624) );
  NAND2X1 U577 ( .A(n1423), .B(N746), .Y(n1080) );
  OAI21X1 U578 ( .A0(n1423), .A1(N746), .B0(n1080), .Y(n1430) );
  NOR2X1 U579 ( .A(n1424), .B(n167), .Y(n1423) );
  NOR2X1 U580 ( .A(n1578), .B(n1577), .Y(n1575) );
  OAI31X1 U581 ( .A0(n1575), .A1(n1557), .A2(n1556), .B0(n1555), .Y(n1589) );
  NOR2X1 U582 ( .A(n2655), .B(n2654), .Y(n2695) );
  NOR2X1 U583 ( .A(next_work_cntr[8]), .B(n2697), .Y(n2732) );
  NOR2X1 U584 ( .A(n969), .B(n1359), .Y(n965) );
  NOR2X1 U585 ( .A(n192), .B(n857), .Y(n851) );
  OAI21X1 U586 ( .A0(n973), .A1(n851), .B0(n864), .Y(n852) );
  NOR2X1 U587 ( .A(n1607), .B(n1649), .Y(n1631) );
  NAND2X1 U588 ( .A(n1663), .B(n1662), .Y(n1664) );
  NOR2BX1 U589 ( .AN(n2826), .B(n2860), .Y(n2862) );
  OAI2BB2X1 U590 ( .B0(n1629), .B1(n1628), .A0N(n1629), .A1N(n1628), .Y(n1662)
         );
  OAI31X1 U591 ( .A0(n1527), .A1(n1526), .A2(n1525), .B0(n1524), .Y(n1544) );
  NOR2X1 U592 ( .A(n2756), .B(n2782), .Y(n2760) );
  NOR2BX1 U593 ( .AN(n1551), .B(n1548), .Y(n1525) );
  AND2X2 U594 ( .A(n2173), .B(n2166), .Y(n2160) );
  OAI21X1 U595 ( .A0(n2166), .A1(n2165), .B0(n2164), .Y(n2170) );
  OAI21X1 U596 ( .A0(n2948), .A1(n2947), .B0(n2946), .Y(n2953) );
  OAI2BB2X1 U597 ( .B0(n2648), .B1(n2157), .A0N(n2648), .A1N(n2157), .Y(n2166)
         );
  NOR3X1 U598 ( .A(n2259), .B(n2266), .C(n2254), .Y(n2263) );
  CLKINVX1 U599 ( .A(n2254), .Y(n2251) );
  NOR2X1 U600 ( .A(n2254), .B(n2253), .Y(n2256) );
  OAI2BB2X1 U601 ( .B0(n2251), .B1(n2253), .A0N(n2251), .A1N(n2253), .Y(n2275)
         );
  OAI2BB2X1 U602 ( .B0(next_work_cntr[7]), .B1(n2150), .A0N(next_work_cntr[7]), 
        .A1N(n2150), .Y(n2254) );
  OAI2BB2X1 U603 ( .B0(n2826), .B1(n2860), .A0N(n2826), .A1N(n2860), .Y(n2880)
         );
  OAI21X1 U604 ( .A0(n1738), .A1(n1737), .B0(n1736), .Y(n1745) );
  NOR2X1 U605 ( .A(N2282), .B(n1859), .Y(n1854) );
  OAI21X1 U606 ( .A0(n1842), .A1(n199), .B0(n1847), .Y(n1859) );
  AOI22X1 U607 ( .A0(n1862), .A1(n1861), .B0(n1860), .B1(n1859), .Y(n2111) );
  NOR2X2 U608 ( .A(n41), .B(n2486), .Y(next_work_cntr[1]) );
  OAI21X1 U609 ( .A0(n194), .A1(n1807), .B0(n1806), .Y(n1812) );
  OAI31X1 U610 ( .A0(n1786), .A1(work_cntr[9]), .A2(n1785), .B0(n1784), .Y(
        n1791) );
  OAI21X1 U611 ( .A0(n160), .A1(n1776), .B0(n1780), .Y(n1785) );
  OAI2BB2X1 U612 ( .B0(n152), .B1(n2326), .A0N(n152), .A1N(n2326), .Y(n2330)
         );
  NOR2X2 U613 ( .A(n161), .B(n1031), .Y(n2326) );
  OAI21X1 U614 ( .A0(n1071), .A1(n1069), .B0(cr_read_cntr[4]), .Y(n1070) );
  OAI31X1 U615 ( .A0(n2494), .A1(n2493), .A2(n2492), .B0(n2491), .Y(n2497) );
  OAI21X1 U616 ( .A0(n2482), .A1(n2481), .B0(n2480), .Y(n2492) );
  AOI221X1 U617 ( .A0(n1287), .A1(n1286), .B0(n1285), .B1(n1286), .C0(n1294), 
        .Y(n1289) );
  OAI21X1 U618 ( .A0(n1007), .A1(n1006), .B0(n1005), .Y(n1285) );
  OAI2BB2X1 U619 ( .B0(work_cntr[6]), .B1(n1242), .A0N(work_cntr[6]), .A1N(
        n1242), .Y(n1252) );
  NAND2X1 U620 ( .A(n2500), .B(n1254), .Y(n1242) );
  OAI2BB2X1 U621 ( .B0(n1222), .B1(n1221), .A0N(n1222), .A1N(n1220), .Y(n1230)
         );
  OAI21X1 U622 ( .A0(n197), .A1(n1823), .B0(n1822), .Y(n1828) );
  OAI21X1 U623 ( .A0(n184), .A1(n1755), .B0(n1754), .Y(n1760) );
  OAI31X1 U624 ( .A0(n1004), .A1(n1003), .A2(n1002), .B0(n1001), .Y(n1295) );
  OAI21X1 U625 ( .A0(n988), .A1(n987), .B0(n986), .Y(n1002) );
  NOR2X1 U626 ( .A(n971), .B(n972), .Y(n981) );
  OAI21X1 U627 ( .A0(n961), .A1(n960), .B0(n959), .Y(n971) );
  OAI21X1 U628 ( .A0(n1468), .A1(n1466), .B0(n1467), .Y(n1516) );
  OAI21X1 U629 ( .A0(n1494), .A1(n1487), .B0(n1466), .Y(n1467) );
  OAI22X2 U630 ( .A0(work_cntr[4]), .A1(n1865), .B0(n164), .B1(n1254), .Y(
        n1267) );
  CLKINVX2 U631 ( .A(n1254), .Y(n1865) );
  CLKINVX1 U632 ( .A(n2099), .Y(n2956) );
  OAI22X1 U633 ( .A0(N2283), .A1(n2099), .B0(n199), .B1(n2956), .Y(n2310) );
  NOR2X1 U634 ( .A(N2282), .B(N205), .Y(n2099) );
  AOI2BB2X2 U635 ( .B0(n1178), .B1(n1181), .A0N(n1178), .A1N(n1177), .Y(n1192)
         );
  OAI21X1 U636 ( .A0(n1171), .A1(n181), .B0(n1170), .Y(n1181) );
  OAI21X1 U637 ( .A0(n2500), .A1(n2600), .B0(n1958), .Y(n2058) );
  NAND2X1 U638 ( .A(n2500), .B(n2600), .Y(n1958) );
  NOR2X1 U639 ( .A(n2047), .B(n2046), .Y(n2050) );
  OAI21X1 U640 ( .A0(n2035), .A1(n193), .B0(n2034), .Y(n2047) );
  NOR2X1 U641 ( .A(n2608), .B(n1966), .Y(n2516) );
  NAND2X1 U642 ( .A(n911), .B(n910), .Y(n916) );
  OAI22X1 U643 ( .A0(n894), .A1(n893), .B0(n897), .B1(n895), .Y(n910) );
  OA21X2 U644 ( .A0(n922), .A1(n921), .B0(n920), .Y(n941) );
  AND2X2 U645 ( .A(n922), .B(n2140), .Y(n924) );
  OAI22X1 U646 ( .A0(n1057), .A1(n1334), .B0(n2135), .B1(n1335), .Y(n922) );
  OAI21X1 U647 ( .A0(n2513), .A1(n2512), .B0(n2511), .Y(n2526) );
  OAI22X1 U648 ( .A0(n161), .A1(n2506), .B0(work_cntr[18]), .B1(n2505), .Y(
        n2512) );
  OAI21X1 U649 ( .A0(n2065), .A1(n2064), .B0(n2063), .Y(n2073) );
  OAI2BB2X1 U650 ( .B0(n1929), .B1(n1928), .A0N(n1929), .A1N(n1927), .Y(n1947)
         );
  OAI22X1 U651 ( .A0(n1917), .A1(n1916), .B0(n1915), .B1(n1914), .Y(n1929) );
  OAI22X1 U652 ( .A0(n1906), .A1(n1914), .B0(n1905), .B1(n1915), .Y(n1928) );
  OAI22X1 U653 ( .A0(n1900), .A1(n1899), .B0(n1901), .B1(n1903), .Y(n1905) );
  OAI21X1 U654 ( .A0(n1645), .A1(n1644), .B0(n1643), .Y(n1668) );
  OAI21X1 U655 ( .A0(n1615), .A1(n1618), .B0(n1613), .Y(n1644) );
  NOR2X1 U656 ( .A(next_work_cntr[15]), .B(next_work_cntr[16]), .Y(n2156) );
  NOR2X4 U657 ( .A(n41), .B(n2353), .Y(next_work_cntr[15]) );
  NOR2X1 U658 ( .A(next_work_cntr[15]), .B(n2672), .Y(n2688) );
  NOR2X1 U659 ( .A(n1378), .B(n1406), .Y(n1434) );
  CLKINVX1 U660 ( .A(n1389), .Y(n63) );
  OAI21X1 U661 ( .A0(n2874), .A1(n2873), .B0(n2872), .Y(n2892) );
  OAI22X1 U662 ( .A0(n2841), .A1(n2840), .B0(n2839), .B1(n2843), .Y(n2874) );
  OAI21X1 U663 ( .A0(n980), .A1(n979), .B0(n978), .Y(n993) );
  AND2X2 U664 ( .A(n980), .B(n2137), .Y(n972) );
  OAI22X1 U665 ( .A0(n1355), .A1(n1133), .B0(n1359), .B1(n2134), .Y(n980) );
  OAI22X1 U666 ( .A0(n1090), .A1(n1089), .B0(n1097), .B1(n1088), .Y(n1116) );
  OAI21X1 U667 ( .A0(n1061), .A1(n1060), .B0(n1059), .Y(n1097) );
  OAI22X1 U668 ( .A0(n1113), .A1(n1112), .B0(n1114), .B1(n1111), .Y(n1131) );
  OAI21X1 U669 ( .A0(n1100), .A1(n1099), .B0(n1098), .Y(n1114) );
  INVXL U670 ( .A(n925), .Y(n64) );
  CLKINVX1 U671 ( .A(n64), .Y(n65) );
  NOR2X1 U672 ( .A(n2695), .B(n2693), .Y(n2685) );
  NOR2X1 U673 ( .A(n2666), .B(n2692), .Y(n2693) );
  NOR2X1 U674 ( .A(n2749), .B(n2747), .Y(n2730) );
  OAI2BB2X1 U675 ( .B0(n1523), .B1(n1522), .A0N(n1523), .A1N(n1522), .Y(n1542)
         );
  AOI211X1 U676 ( .A0(n354), .A1(n1317), .B0(n1158), .C0(n1159), .Y(n711) );
  OAI31X1 U677 ( .A0(n255), .A1(n1329), .A2(n1328), .B0(n1327), .Y(n1336) );
  AOI211X4 U678 ( .A0(n1333), .A1(n1334), .B0(n1332), .C0(n1331), .Y(n1338) );
  OAI31X1 U679 ( .A0(n255), .A1(n1325), .A2(n1324), .B0(n1323), .Y(n1333) );
  CLKINVX1 U680 ( .A(n1513), .Y(n66) );
  CLKINVX1 U681 ( .A(n66), .Y(n67) );
  OAI31X1 U682 ( .A0(n1633), .A1(n1621), .A2(n1620), .B0(n1619), .Y(n1636) );
  NOR2X1 U683 ( .A(n929), .B(n937), .Y(n940) );
  CLKINVX1 U684 ( .A(n2149), .Y(n68) );
  CLKINVX1 U685 ( .A(n2933), .Y(n69) );
  NAND3X1 U686 ( .A(work_cntr[4]), .B(work_cntr[5]), .C(n68), .Y(n1045) );
  NOR2X1 U687 ( .A(n1193), .B(n1192), .Y(n1197) );
  AOI2BB2X2 U688 ( .B0(n1189), .B1(n1188), .A0N(n1189), .A1N(n1193), .Y(n1199)
         );
  AOI2BB2X2 U689 ( .B0(work_cntr[15]), .B1(n1186), .A0N(n1176), .A1N(n1201), 
        .Y(n1193) );
  NAND2X1 U690 ( .A(n2014), .B(n1863), .Y(n1966) );
  NAND2X1 U691 ( .A(n181), .B(n1863), .Y(n1444) );
  NOR4X2 U692 ( .A(work_cntr[13]), .B(work_cntr[15]), .C(n256), .D(n1438), .Y(
        n1863) );
  NOR2BX1 U693 ( .AN(n451), .B(curr_time[2]), .Y(n377) );
  AOI31X1 U694 ( .A0(n1028), .A1(curr_time[2]), .A2(n376), .B0(n377), .Y(n428)
         );
  OAI211X1 U695 ( .A0(curr_time[2]), .A1(n1028), .B0(curr_time[1]), .C0(n1030), 
        .Y(n374) );
  CLKINVX1 U696 ( .A(n723), .Y(\im_a[1]_BAR ) );
  CLKINVX1 U697 ( .A(n725), .Y(\im_a[2]_BAR ) );
  CLKINVX1 U698 ( .A(n727), .Y(\im_a[3]_BAR ) );
  CLKINVX1 U699 ( .A(n729), .Y(\im_a[4]_BAR ) );
  CLKINVX1 U700 ( .A(n731), .Y(\im_a[5]_BAR ) );
  CLKINVX1 U701 ( .A(n733), .Y(\im_a[6]_BAR ) );
  CLKINVX1 U702 ( .A(n735), .Y(\im_a[7]_BAR ) );
  CLKINVX1 U703 ( .A(n737), .Y(\im_a[8]_BAR ) );
  CLKINVX1 U704 ( .A(n739), .Y(\im_a[9]_BAR ) );
  CLKINVX1 U705 ( .A(n741), .Y(\im_a[10]_BAR ) );
  CLKINVX1 U706 ( .A(n743), .Y(\im_a[11]_BAR ) );
  CLKINVX1 U707 ( .A(n745), .Y(\im_a[12]_BAR ) );
  CLKINVX1 U708 ( .A(n747), .Y(\im_a[13]_BAR ) );
  CLKINVX1 U709 ( .A(n749), .Y(\im_a[14]_BAR ) );
  CLKINVX1 U710 ( .A(n751), .Y(\im_a[15]_BAR ) );
  CLKINVX1 U711 ( .A(n753), .Y(\im_a[16]_BAR ) );
  CLKINVX1 U712 ( .A(n755), .Y(\im_a[17]_BAR ) );
  CLKINVX1 U713 ( .A(n758), .Y(\im_a[18]_BAR ) );
  NOR3X2 U714 ( .A(n468), .B(n467), .C(n466), .Y(\DP_OP_280J1_126_7605/I2 ) );
  CLKINVX1 U715 ( .A(n409), .Y(n468) );
  NAND2X1 U716 ( .A(n1907), .B(n1949), .Y(n1912) );
  NAND2X1 U717 ( .A(write_cntr[6]), .B(n1949), .Y(n1924) );
  NOR2X1 U718 ( .A(n1949), .B(n363), .Y(n381) );
  AOI211X4 U719 ( .A0(\intadd_3/SUM[7] ), .A1(n251), .B0(n1365), .C0(n339), 
        .Y(n659) );
  OAI21X1 U720 ( .A0(write_addr[10]), .A1(n1313), .B0(n1312), .Y(n1315) );
  OAI2BB2X1 U721 ( .B0(n1312), .B1(n153), .A0N(n1312), .A1N(n153), .Y(n1364)
         );
  NOR2X1 U722 ( .A(n1312), .B(n153), .Y(n1073) );
  NAND2X1 U723 ( .A(n1713), .B(n1367), .Y(n1312) );
  CLKINVX1 U724 ( .A(next_work_cntr[18]), .Y(n2648) );
  NOR2X2 U725 ( .A(n41), .B(n2329), .Y(next_work_cntr[18]) );
  OAI211X1 U726 ( .A0(n1455), .A1(n1454), .B0(n1453), .C0(n1452), .Y(n1466) );
  NAND4X1 U727 ( .A(n1449), .B(n1465), .C(n1456), .D(n1443), .Y(n1454) );
  NOR2X1 U728 ( .A(write_cntr[8]), .B(n1951), .Y(n1893) );
  NAND2X1 U729 ( .A(n1880), .B(n1951), .Y(n1886) );
  NAND2X1 U730 ( .A(n1951), .B(write_cntr[8]), .Y(n1892) );
  OAI31X1 U731 ( .A0(n1241), .A1(n1240), .A2(n1239), .B0(n1238), .Y(n1247) );
  OAI2BB2X2 U732 ( .B0(work_cntr[8]), .B1(n1227), .A0N(work_cntr[8]), .A1N(
        n1227), .Y(n1241) );
  OAI21X1 U733 ( .A0(n416), .A1(n415), .B0(n452), .Y(n460) );
  NAND2X1 U734 ( .A(n414), .B(n413), .Y(n452) );
  OAI21X1 U735 ( .A0(n397), .A1(n396), .B0(n434), .Y(n458) );
  OA21X1 U736 ( .A0(m_1[2]), .A1(n1019), .B0(n1020), .Y(n397) );
  AOI2BB2X2 U737 ( .B0(n1499), .B1(n1498), .A0N(n1499), .A1N(n1498), .Y(n1578)
         );
  NOR2BX1 U738 ( .AN(n1499), .B(n1498), .Y(n1531) );
  OAI2BB2X2 U739 ( .B0(n1479), .B1(n1478), .A0N(n1479), .A1N(n1478), .Y(n1499)
         );
  INVXL U740 ( .A(n698), .Y(n70) );
  CLKINVX1 U741 ( .A(n70), .Y(n71) );
  OAI22X2 U742 ( .A0(n2548), .A1(n2547), .B0(work_cntr[12]), .B1(n2546), .Y(
        n2565) );
  CLKINVX1 U743 ( .A(n2547), .Y(n2546) );
  NOR2X2 U744 ( .A(n234), .B(n1391), .Y(n1397) );
  NOR2X1 U745 ( .A(n1717), .B(n508), .Y(n551) );
  NOR2X1 U746 ( .A(n235), .B(n1717), .Y(n1716) );
  NAND2BX1 U747 ( .AN(n1715), .B(n770), .Y(n1717) );
  NOR2X1 U748 ( .A(n1402), .B(n352), .Y(n632) );
  CLKINVX1 U749 ( .A(n348), .Y(n640) );
  NAND2BX1 U750 ( .AN(n1393), .B(n347), .Y(n348) );
  AOI211X4 U751 ( .A0(\intadd_3/SUM[5] ), .A1(n251), .B0(n1371), .C0(n327), 
        .Y(n668) );
  AOI211X4 U752 ( .A0(n179), .A1(n251), .B0(n1382), .C0(n342), .Y(n648) );
  OAI21X2 U753 ( .A0(n1429), .A1(n1428), .B0(n333), .Y(n692) );
  OAI211X1 U754 ( .A0(n457), .A1(n474), .B0(n456), .C0(n455), .Y(\C1/Z_1 ) );
  OAI211X1 U755 ( .A0(n422), .A1(n474), .B0(n421), .C0(n420), .Y(\C1/Z_3 ) );
  NAND2X1 U756 ( .A(n468), .B(n408), .Y(n474) );
  NOR2X1 U757 ( .A(n1612), .B(n1611), .Y(n1594) );
  CLKINVX1 U758 ( .A(n1589), .Y(n1612) );
  NAND2X1 U759 ( .A(n1603), .B(n1590), .Y(n1618) );
  NOR3X1 U760 ( .A(n1607), .B(n1641), .C(n1608), .Y(n1603) );
  NOR2X1 U761 ( .A(n2600), .B(n1045), .Y(n1044) );
  OAI21X2 U762 ( .A0(n256), .A1(n1036), .B0(n1035), .Y(n2356) );
  NAND2X1 U763 ( .A(n256), .B(n1036), .Y(n1035) );
  AOI222X4 U764 ( .A0(n4), .A1(n777), .B0(n776), .B1(n102), .C0(n251), .C1(
        \intadd_3/SUM[8] ), .Y(n654) );
  NAND2BX1 U765 ( .AN(n1627), .B(n1626), .Y(n1660) );
  CLKINVX1 U766 ( .A(n2153), .Y(next_work_cntr[14]) );
  NAND2X1 U767 ( .A(n257), .B(n2360), .Y(n2153) );
  OAI21X1 U768 ( .A0(n2545), .A1(n2544), .B0(n2543), .Y(n2552) );
  OAI22X1 U769 ( .A0(n2545), .A1(n2536), .B0(n2535), .B1(n2534), .Y(n2540) );
  CLKINVX1 U770 ( .A(n2538), .Y(n2545) );
  NOR4X1 U771 ( .A(next_work_cntr[9]), .B(n2656), .C(n2680), .D(n2691), .Y(
        n2666) );
  NOR2X1 U772 ( .A(n2680), .B(n2679), .Y(n2715) );
  NAND2BX1 U773 ( .AN(next_work_cntr[13]), .B(n2650), .Y(n2680) );
  OAI21X2 U774 ( .A0(n371), .A1(n370), .B0(n369), .Y(n376) );
  NOR2X1 U775 ( .A(work_cntr[17]), .B(n2515), .Y(n2506) );
  OAI21X2 U776 ( .A0(n2516), .A1(n181), .B0(n2515), .Y(n2525) );
  NAND2X1 U777 ( .A(n2516), .B(n181), .Y(n2515) );
  AND2X2 U778 ( .A(n350), .B(n349), .Y(n636) );
  CLKINVX1 U779 ( .A(n2661), .Y(next_work_cntr[16]) );
  OAI21X2 U780 ( .A0(n2159), .A1(n2661), .B0(n2158), .Y(n2162) );
  NAND2X1 U781 ( .A(n257), .B(n2337), .Y(n2661) );
  OAI2BB2X1 U782 ( .B0(next_work_cntr[13]), .B1(n2193), .A0N(
        next_work_cntr[13]), .A1N(n2193), .Y(n2191) );
  NOR2X1 U783 ( .A(next_work_cntr[13]), .B(n2193), .Y(n2154) );
  NAND2X1 U784 ( .A(n2152), .B(n2650), .Y(n2193) );
  NOR2X1 U785 ( .A(n2629), .B(n2628), .Y(n2630) );
  NOR2X2 U786 ( .A(N2283), .B(N2282), .Y(n2628) );
  AOI211X4 U787 ( .A0(\intadd_3/SUM[6] ), .A1(n251), .B0(n1316), .C0(n324), 
        .Y(n664) );
  CLKINVX1 U788 ( .A(n2453), .Y(n2457) );
  OAI22X1 U789 ( .A0(work_cntr[4]), .A1(n68), .B0(n164), .B1(n2149), .Y(n2453)
         );
  AOI2BB2X2 U790 ( .B0(n2786), .B1(n2785), .A0N(n2786), .A1N(n2785), .Y(n2836)
         );
  CLKINVX1 U791 ( .A(n2723), .Y(n2786) );
  OAI211X4 U792 ( .A0(n1304), .A1(n1107), .B0(n1106), .C0(n1105), .Y(n1125) );
  OAI31X4 U793 ( .A0(n2075), .A1(n2072), .A2(n2071), .B0(n2070), .Y(n2076) );
  OAI21X2 U794 ( .A0(n1165), .A1(n1428), .B0(n1164), .Y(n2145) );
  CLKINVX1 U795 ( .A(n1497), .Y(n1533) );
  OAI2BB2X1 U796 ( .B0(n2548), .B1(n1463), .A0N(n2548), .A1N(n1463), .Y(n1497)
         );
  AOI22X1 U797 ( .A0(n1210), .A1(n1209), .B0(n1208), .B1(n1216), .Y(n1219) );
  OAI21X2 U798 ( .A0(n1203), .A1(n2548), .B0(n1202), .Y(n1216) );
  OAI31X1 U799 ( .A0(n2291), .A1(n2290), .A2(n2289), .B0(n2288), .Y(n2302) );
  AOI211X4 U800 ( .A0(n2278), .A1(n2277), .B0(work_cntr[4]), .C0(n41), .Y(
        n2291) );
  CLKINVX1 U801 ( .A(n72), .Y(n73) );
  AND2X2 U802 ( .A(n345), .B(n344), .Y(n644) );
  CLKINVX1 U803 ( .A(n74), .Y(n75) );
  NOR2X2 U804 ( .A(N2284), .B(n2082), .Y(n2102) );
  OAI21X1 U805 ( .A0(n2784), .A1(n2797), .B0(n80), .Y(n2785) );
  NAND2X1 U806 ( .A(n2778), .B(n2797), .Y(n2812) );
  NOR2BX2 U807 ( .AN(n2773), .B(n2822), .Y(n2797) );
  NAND2X1 U808 ( .A(n1896), .B(n1950), .Y(n1897) );
  CLKINVX1 U809 ( .A(n2184), .Y(n76) );
  NAND2X1 U810 ( .A(n1673), .B(n1672), .Y(n1686) );
  NAND2X2 U811 ( .A(n257), .B(n2402), .Y(n2686) );
  CLKINVX1 U812 ( .A(n2402), .Y(n2410) );
  AOI21X2 U813 ( .A0(n187), .A1(n1041), .B0(n1040), .Y(n2402) );
  OAI21X2 U814 ( .A0(n2561), .A1(n187), .B0(n2560), .Y(n2582) );
  NAND2X1 U815 ( .A(n2561), .B(n187), .Y(n2560) );
  NOR2X1 U816 ( .A(work_cntr[8]), .B(n2575), .Y(n2561) );
  CLKINVX1 U817 ( .A(n609), .Y(n618) );
  CLKINVX1 U818 ( .A(n2728), .Y(n77) );
  NOR3BX1 U819 ( .AN(n2886), .B(next_work_cntr[0]), .C(n2885), .Y(n2905) );
  CLKINVX1 U820 ( .A(n2897), .Y(next_work_cntr[0]) );
  OAI21X1 U821 ( .A0(n2607), .A1(n2606), .B0(n2605), .Y(n2614) );
  OAI2BB2X2 U822 ( .B0(work_cntr[6]), .B1(n2591), .A0N(work_cntr[6]), .A1N(
        n2591), .Y(n2606) );
  OAI21X1 U823 ( .A0(n1725), .A1(n1731), .B0(n1724), .Y(n1727) );
  NAND2X1 U824 ( .A(n1960), .B(n1731), .Y(n1455) );
  NOR2X2 U825 ( .A(n152), .B(n1445), .Y(n1731) );
  OAI21X1 U826 ( .A0(n1404), .A1(n207), .B0(n257), .Y(n1317) );
  OAI211X4 U827 ( .A0(n1410), .A1(n1082), .B0(n774), .C0(n1081), .Y(n1404) );
  CLKINVX1 U828 ( .A(n997), .Y(n2132) );
  OAI21X1 U829 ( .A0(n864), .A1(n201), .B0(n863), .Y(n997) );
  CLKINVX1 U830 ( .A(n2753), .Y(n78) );
  OAI21X2 U831 ( .A0(n2576), .A1(n194), .B0(n2575), .Y(n2597) );
  NAND2X1 U832 ( .A(n2576), .B(n194), .Y(n2575) );
  OAI22X2 U833 ( .A0(write_cntr[0]), .A1(n973), .B0(n203), .B1(n864), .Y(n1160) );
  NAND3X1 U834 ( .A(N743), .B(N742), .C(N744), .Y(n1424) );
  OAI21X1 U835 ( .A0(n1995), .A1(n184), .B0(n1959), .Y(n1997) );
  NAND2X1 U836 ( .A(n1995), .B(n184), .Y(n1959) );
  NOR2X2 U837 ( .A(n1175), .B(n1438), .Y(n1995) );
  CLKINVX1 U838 ( .A(n2807), .Y(n2830) );
  NAND2X1 U839 ( .A(n2609), .B(n2500), .Y(n2591) );
  OAI22X2 U840 ( .A0(n2609), .A1(n164), .B0(n2608), .B1(work_cntr[4]), .Y(
        n2626) );
  NOR2X2 U841 ( .A(n2629), .B(N2284), .Y(n2609) );
  CLKINVX1 U842 ( .A(n1276), .Y(n1278) );
  OAI21X1 U843 ( .A0(n1273), .A1(n2462), .B0(n1272), .Y(n1276) );
  CLKINVX1 U844 ( .A(n2654), .Y(next_work_cntr[19]) );
  NAND2X1 U845 ( .A(n257), .B(n2330), .Y(n2654) );
  OAI2BB2X2 U846 ( .B0(next_work_cntr[8]), .B1(n2697), .A0N(next_work_cntr[8]), 
        .A1N(n2697), .Y(n2749) );
  NOR2BX1 U847 ( .AN(n2717), .B(n2719), .Y(n2697) );
  INVXL U848 ( .A(n2783), .Y(n79) );
  CLKINVX1 U849 ( .A(n79), .Y(n80) );
  CLKINVX1 U850 ( .A(n2684), .Y(next_work_cntr[11]) );
  NAND2X1 U851 ( .A(n257), .B(n2384), .Y(n2684) );
  INVXL U852 ( .A(n1529), .Y(n81) );
  CLKINVX1 U853 ( .A(n81), .Y(n82) );
  OAI2BB2X1 U854 ( .B0(n1319), .B1(n2133), .A0N(n1319), .A1N(n2133), .Y(n999)
         );
  NOR2BX2 U855 ( .AN(n2133), .B(n989), .Y(n994) );
  OAI31X4 U856 ( .A0(n2039), .A1(n2032), .A2(n2031), .B0(n2030), .Y(n2036) );
  NOR2BX2 U857 ( .AN(n2016), .B(n2013), .Y(n2039) );
  OAI21X1 U858 ( .A0(n1477), .A1(n2501), .B0(n1462), .Y(n1463) );
  NAND2BX1 U859 ( .AN(n2501), .B(n2548), .Y(n1438) );
  OAI22X1 U860 ( .A0(n2501), .A1(n1201), .B0(n1196), .B1(n180), .Y(n1212) );
  NOR2X1 U861 ( .A(n2501), .B(n2560), .Y(n2547) );
  NAND2X1 U862 ( .A(n160), .B(n180), .Y(n2501) );
  OAI21X2 U863 ( .A0(work_cntr[12]), .A1(n1038), .B0(n1037), .Y(n2375) );
  NAND2X1 U864 ( .A(work_cntr[12]), .B(n1038), .Y(n1037) );
  NOR2X1 U865 ( .A(n180), .B(n1039), .Y(n1038) );
  ADDFX2 U866 ( .A(n1297), .B(n1291), .CI(n1290), .CO(n1412), .S(n1165) );
  NOR2X1 U867 ( .A(n1298), .B(n1297), .Y(n1303) );
  CLKINVX1 U868 ( .A(n1299), .Y(n1297) );
  NOR2BX1 U869 ( .AN(n1320), .B(n1325), .Y(n1329) );
  CLKINVX1 U870 ( .A(n1321), .Y(n1320) );
  OAI22X1 U871 ( .A0(n976), .A1(n1361), .B0(n2137), .B1(n1375), .Y(n989) );
  CLKINVX1 U872 ( .A(n1375), .Y(n1361) );
  NOR2X2 U873 ( .A(n409), .B(n408), .Y(n473) );
  AND2X2 U874 ( .A(n467), .B(n366), .Y(n472) );
  OAI2BB2X2 U875 ( .B0(n2271), .B1(n2270), .A0N(n2271), .A1N(n2270), .Y(n2290)
         );
  AOI2BB2X2 U876 ( .B0(work_cntr[10]), .B1(n1477), .A0N(work_cntr[10]), .A1N(
        n1477), .Y(n1479) );
  NOR2X1 U877 ( .A(n1438), .B(n1477), .Y(n1441) );
  NAND2X2 U878 ( .A(work_cntr[19]), .B(n1437), .Y(n1477) );
  CLKINVX1 U879 ( .A(n856), .Y(n2143) );
  AOI2BB2X2 U880 ( .B0(n856), .B1(n855), .A0N(n856), .A1N(n855), .Y(n1056) );
  NAND3X1 U881 ( .A(n891), .B(n856), .C(n881), .Y(n859) );
  OAI22X2 U882 ( .A0(n864), .A1(n189), .B0(n973), .B1(n850), .Y(n856) );
  INVXL U883 ( .A(n964), .Y(n83) );
  CLKINVX1 U884 ( .A(n83), .Y(n84) );
  NAND2X1 U885 ( .A(n2733), .B(n2734), .Y(n2747) );
  NAND2X2 U886 ( .A(n257), .B(n2422), .Y(n2733) );
  OAI21X1 U887 ( .A0(n2450), .A1(n2449), .B0(n2448), .Y(n2456) );
  OAI21X1 U888 ( .A0(n2300), .A1(n2299), .B0(n2298), .Y(n2307) );
  NOR2X1 U889 ( .A(n2299), .B(n2300), .Y(n2289) );
  NAND2X1 U890 ( .A(n2287), .B(n2286), .Y(n2300) );
  AOI222X4 U891 ( .A0(\intadd_3/SUM[3] ), .A1(n251), .B0(n776), .B1(N748), 
        .C0(n774), .C1(n1434), .Y(n677) );
  CLKINVX1 U892 ( .A(n1355), .Y(n1359) );
  NAND2X1 U893 ( .A(n956), .B(n958), .Y(n1355) );
  CLKINVX1 U894 ( .A(n866), .Y(n874) );
  OAI22X1 U895 ( .A0(n2068), .A1(n2073), .B0(n2148), .B1(n2067), .Y(n2085) );
  NOR2X1 U896 ( .A(n2148), .B(n2073), .Y(n2081) );
  OAI22X2 U897 ( .A0(work_cntr[4]), .A1(n197), .B0(n164), .B1(work_cntr[5]), 
        .Y(n2148) );
  CLKINVX1 U898 ( .A(n2139), .Y(n1119) );
  OAI2BB1X2 U899 ( .A0N(n191), .A1N(n865), .B0(n906), .Y(n2139) );
  AOI221X4 U900 ( .A0(n2652), .A1(next_work_cntr[14]), .B0(n2669), .B1(
        next_work_cntr[14]), .C0(n2675), .Y(n2714) );
  NOR2X2 U901 ( .A(n2651), .B(n2653), .Y(n2675) );
  CLKINVX1 U902 ( .A(n868), .Y(n867) );
  OAI21X2 U903 ( .A0(work_cntr[8]), .A1(n1042), .B0(n1041), .Y(n2413) );
  NAND2X1 U904 ( .A(work_cntr[8]), .B(n1042), .Y(n1041) );
  CLKINVX1 U905 ( .A(n1043), .Y(n1042) );
  OAI21X2 U906 ( .A0(n1962), .A1(n152), .B0(n2955), .Y(n1979) );
  NOR2X2 U907 ( .A(n1175), .B(n1437), .Y(n1962) );
  CLKINVX1 U908 ( .A(n2322), .Y(n781) );
  CLKINVX1 U909 ( .A(\DP_OP_280J1_126_7605/I3 ), .Y(n85) );
  NAND2X1 U910 ( .A(n257), .B(n2148), .Y(n2271) );
  NAND2X1 U911 ( .A(n146), .B(n257), .Y(n2897) );
  NAND3X1 U912 ( .A(n2149), .B(n1865), .C(n257), .Y(n2820) );
  OAI21X1 U913 ( .A0(n1433), .A1(n712), .B0(n713), .Y(n628) );
  OAI21X1 U914 ( .A0(n1433), .A1(n136), .B0(n2147), .Y(n683) );
  OA21X2 U915 ( .A0(n1433), .A1(n213), .B0(n2146), .Y(n685) );
  NOR2X1 U916 ( .A(n612), .B(n1433), .Y(n553) );
  OAI222X4 U917 ( .A0(n211), .A1(n1433), .B0(n1431), .B1(n1422), .C0(n1428), 
        .C1(n1421), .Y(n696) );
  CLKINVX1 U918 ( .A(n776), .Y(n1433) );
  INVXL U919 ( .A(n1685), .Y(n86) );
  CLKINVX1 U920 ( .A(n86), .Y(n87) );
  OAI22X2 U921 ( .A0(write_cntr[3]), .A1(n957), .B0(n200), .B1(n975), .Y(n2137) );
  NOR2X1 U922 ( .A(n973), .B(n931), .Y(n957) );
  CLKINVX1 U923 ( .A(n2462), .Y(n2470) );
  NOR2X1 U924 ( .A(n68), .B(n1254), .Y(n2462) );
  CLKINVX1 U925 ( .A(n1057), .Y(n2135) );
  OAI22X2 U926 ( .A0(n195), .A1(n864), .B0(n973), .B1(n858), .Y(n1057) );
  OAI22X2 U927 ( .A0(n1101), .A1(n1298), .B0(n2140), .B1(n1308), .Y(n1123) );
  CLKINVX1 U928 ( .A(n2140), .Y(n1101) );
  CLKINVX1 U929 ( .A(n2384), .Y(n2671) );
  AOI21X1 U930 ( .A0(n180), .A1(n1039), .B0(n1038), .Y(n2384) );
  AND2X2 U931 ( .A(write_addr[15]), .B(n88), .Y(n773) );
  OAI21X1 U932 ( .A0(write_addr[15]), .A1(n1390), .B0(n1389), .Y(n1392) );
  NAND3X2 U933 ( .A(n718), .B(n717), .C(n2969), .Y(n760) );
  NAND2X1 U934 ( .A(n598), .B(n597), .Y(n609) );
  OAI21X1 U935 ( .A0(n1714), .A1(n597), .B0(n598), .Y(n581) );
  OAI21X1 U936 ( .A0(n551), .A1(n597), .B0(n598), .Y(n562) );
  OA21X2 U937 ( .A0(n514), .A1(n513), .B0(n1696), .Y(n598) );
  NAND2X2 U938 ( .A(n1115), .B(n1114), .Y(n1305) );
  NOR2X1 U939 ( .A(n869), .B(n871), .Y(n872) );
  OAI22X2 U940 ( .A0(n160), .A1(n1218), .B0(n2541), .B1(n1865), .Y(n1229) );
  OAI21X2 U941 ( .A0(n2014), .A1(n160), .B0(n2541), .Y(n2026) );
  NAND2X2 U942 ( .A(n2014), .B(n160), .Y(n2541) );
  NAND2X1 U943 ( .A(n891), .B(next_cr_x[6]), .Y(n1051) );
  OAI21X2 U944 ( .A0(n891), .A1(next_cr_x[6]), .B0(n1051), .Y(n1093) );
  AOI221X4 U945 ( .A0(n854), .A1(n192), .B0(n865), .B1(n192), .C0(n853), .Y(
        n891) );
  INVX3 U946 ( .A(n2482), .Y(n2476) );
  OAI22X2 U947 ( .A0(N2283), .A1(n2120), .B0(n199), .B1(n1047), .Y(n2482) );
  NOR2X1 U948 ( .A(n153), .B(n1363), .Y(n1379) );
  NOR2X2 U949 ( .A(n1720), .B(n153), .Y(n770) );
  OAI21X1 U950 ( .A0(n1076), .A1(write_addr[18]), .B0(n1083), .Y(n1403) );
  INVX3 U951 ( .A(n718), .Y(n716) );
  AOI21X1 U952 ( .A0(n184), .A1(n1037), .B0(n1036), .Y(n2652) );
  NOR2X2 U953 ( .A(read_cntr[0]), .B(read_cntr[1]), .Y(n619) );
  NAND2X1 U954 ( .A(read_cntr[0]), .B(n172), .Y(n1869) );
  NOR2X1 U955 ( .A(read_cntr[0]), .B(n719), .Y(n670) );
  NAND2X1 U956 ( .A(n63), .B(write_addr[16]), .Y(n1077) );
  NAND2X1 U957 ( .A(n2014), .B(n1254), .Y(n1201) );
  NAND2X1 U958 ( .A(n1254), .B(n1995), .Y(n1202) );
  NOR2X4 U959 ( .A(N2284), .B(n1046), .Y(n1254) );
  INVX16 U960 ( .A(n7), .Y(cr_a[1]) );
  INVX4 U961 ( .A(n779), .Y(n756) );
  INVX16 U962 ( .A(n8), .Y(cr_a[2]) );
  INVX16 U963 ( .A(n5), .Y(cr_a[0]) );
  CLKINVX1 U964 ( .A(n2977), .Y(n93) );
  INVX16 U965 ( .A(n93), .Y(cr_a[3]) );
  CLKINVX1 U966 ( .A(n2975), .Y(n95) );
  INVX16 U967 ( .A(n95), .Y(cr_a[5]) );
  CLKINVX1 U968 ( .A(n2974), .Y(n97) );
  INVX16 U969 ( .A(n97), .Y(cr_a[6]) );
  CLKINVX1 U970 ( .A(n2973), .Y(n99) );
  INVX16 U971 ( .A(n99), .Y(cr_a[7]) );
  INVX16 U972 ( .A(n10), .Y(cr_a[8]) );
  NAND2X1 U973 ( .A(n162), .B(n1604), .Y(n1626) );
  NOR2X1 U974 ( .A(n162), .B(n1604), .Y(n1627) );
  OAI21X1 U975 ( .A0(n162), .A1(n1839), .B0(n1838), .Y(n1844) );
  INVX3 U976 ( .A(n649), .Y(n704) );
  AND2X2 U977 ( .A(n669), .B(n623), .Y(n649) );
  INVX4 U978 ( .A(n715), .Y(n103) );
  NAND2BX1 U979 ( .AN(n1788), .B(n1790), .Y(n1794) );
  NOR2X1 U980 ( .A(n1782), .B(n1787), .Y(n1788) );
  NOR2X1 U981 ( .A(n1287), .B(n1286), .Y(n1284) );
  NOR2X1 U982 ( .A(n1160), .B(n1163), .Y(n1287) );
  NAND2X1 U983 ( .A(n2514), .B(n2524), .Y(n2523) );
  NOR2X1 U984 ( .A(n1546), .B(n1545), .Y(n1553) );
  NAND2X1 U985 ( .A(n2896), .B(n2901), .Y(n2913) );
  NAND2X1 U986 ( .A(n2795), .B(n2805), .Y(n2859) );
  NAND2X1 U987 ( .A(n2816), .B(n2815), .Y(n2805) );
  NOR2BX1 U988 ( .AN(\h_1[2] ), .B(curr_time[19]), .Y(n1012) );
  OAI21X1 U989 ( .A0(n1506), .A1(n1505), .B0(n1504), .Y(n1507) );
  NOR2X2 U990 ( .A(n1484), .B(n1506), .Y(n1526) );
  NOR2X1 U991 ( .A(n193), .B(n1488), .Y(n1506) );
  NOR2BX1 U992 ( .AN(n1579), .B(n1578), .Y(n1530) );
  NOR2X1 U993 ( .A(n1528), .B(n82), .Y(n1579) );
  CLKINVX1 U994 ( .A(n2624), .Y(n2635) );
  AOI21X1 U995 ( .A0(n2624), .A1(n2623), .B0(n2622), .Y(n2638) );
  NOR2BX1 U996 ( .AN(n1592), .B(n1591), .Y(n1561) );
  NAND2X1 U997 ( .A(n1559), .B(n1558), .Y(n1591) );
  OAI21X1 U998 ( .A0(n1788), .A1(n1783), .B0(n187), .Y(n1789) );
  NOR2BX1 U999 ( .AN(n1776), .B(n1775), .Y(n1783) );
  NOR2X1 U1000 ( .A(n2651), .B(n2656), .Y(n2657) );
  NAND2X1 U1001 ( .A(n2156), .B(n2664), .Y(n2656) );
  NOR2X1 U1002 ( .A(n948), .B(n947), .Y(n953) );
  NAND2X1 U1003 ( .A(n2271), .B(n2270), .Y(n2280) );
  OAI21X1 U1004 ( .A0(n2269), .A1(n2268), .B0(n2267), .Y(n2270) );
  AOI211X1 U1005 ( .A0(n1946), .A1(n1945), .B0(n1944), .C0(n1943), .Y(n2129)
         );
  NOR2BX1 U1006 ( .AN(n1932), .B(n1948), .Y(n1946) );
  NAND2X1 U1007 ( .A(n1472), .B(n1484), .Y(n1476) );
  NOR2X1 U1008 ( .A(n1458), .B(n1483), .Y(n1472) );
  NOR2X1 U1009 ( .A(next_work_cntr[8]), .B(n2234), .Y(n2151) );
  NAND2X1 U1010 ( .A(n2150), .B(n2733), .Y(n2234) );
  NOR2BX1 U1011 ( .AN(n2248), .B(n2259), .Y(n2257) );
  NOR2X1 U1012 ( .A(n1976), .B(n1975), .Y(n1984) );
  NOR2X1 U1013 ( .A(n2891), .B(n2889), .Y(n2834) );
  OAI211X4 U1014 ( .A0(n2825), .A1(n2832), .B0(n2824), .C0(n2837), .Y(n2891)
         );
  AOI2BB2X2 U1015 ( .B0(write_cntr[11]), .B1(n1875), .A0N(write_cntr[11]), 
        .A1N(n1875), .Y(n1887) );
  NOR2X1 U1016 ( .A(n204), .B(n1883), .Y(n1875) );
  CLKINVX1 U1017 ( .A(next_work_cntr[8]), .Y(n2690) );
  NOR2X2 U1018 ( .A(n41), .B(n2413), .Y(next_work_cntr[8]) );
  NOR2BX1 U1019 ( .AN(n1244), .B(n1246), .Y(n1249) );
  NOR2X1 U1020 ( .A(n2608), .B(n2541), .Y(n2559) );
  CLKINVX1 U1021 ( .A(n2609), .Y(n2608) );
  NOR2XL U1022 ( .A(n2968), .B(n2967), .Y(n105) );
  CLKINVX1 U1023 ( .A(n2970), .Y(n106) );
  NAND2X1 U1024 ( .A(n669), .B(n2645), .Y(n2967) );
  NOR2BX1 U1025 ( .AN(n1094), .B(n1298), .Y(n1095) );
  NAND2BX1 U1026 ( .AN(n1093), .B(n1091), .Y(n1094) );
  OAI211X1 U1027 ( .A0(n1408), .A1(n1407), .B0(n777), .C0(n1409), .Y(n2944) );
  NAND3X1 U1028 ( .A(n1408), .B(n1406), .C(n1405), .Y(n1409) );
  OAI21X1 U1029 ( .A0(n2846), .A1(n2845), .B0(n2844), .Y(n2873) );
  NAND3X1 U1030 ( .A(write_cntr[8]), .B(write_cntr[7]), .C(n907), .Y(n857) );
  NOR3X2 U1031 ( .A(n191), .B(n931), .C(n841), .Y(n907) );
  NOR2X1 U1032 ( .A(N2283), .B(n2956), .Y(n2107) );
  OAI2BB2X1 U1033 ( .B0(n2599), .B1(n2598), .A0N(n2599), .A1N(n2597), .Y(n2607) );
  OAI21X1 U1034 ( .A0(n2595), .A1(n2594), .B0(n2593), .Y(n2599) );
  NOR2BX1 U1035 ( .AN(n1667), .B(n1648), .Y(n1647) );
  AOI21X1 U1036 ( .A0(n1648), .A1(n1668), .B0(n1647), .Y(n1674) );
  OAI2BB2X1 U1037 ( .B0(n1641), .B1(n1640), .A0N(n1641), .A1N(n1640), .Y(n1648) );
  AOI21X1 U1038 ( .A0(n2096), .A1(n165), .B0(n2103), .Y(n2115) );
  NOR2X1 U1039 ( .A(n2096), .B(n165), .Y(n2103) );
  CLKINVX1 U1040 ( .A(n1633), .Y(n1625) );
  OAI2BB2X2 U1041 ( .B0(n1552), .B1(n1553), .A0N(n1552), .A1N(n1553), .Y(n1633) );
  OAI2BB2X1 U1042 ( .B0(n1207), .B1(n1206), .A0N(n1207), .A1N(n1205), .Y(n1217) );
  OAI21X1 U1043 ( .A0(n1200), .A1(n1199), .B0(n1198), .Y(n1207) );
  NAND2X1 U1044 ( .A(n2714), .B(n2713), .Y(n2702) );
  NOR2BX1 U1045 ( .AN(n2729), .B(n77), .Y(n2713) );
  OAI21X1 U1046 ( .A0(n1653), .A1(n1652), .B0(n1661), .Y(n1655) );
  OAI22X1 U1047 ( .A0(n2603), .A1(n2606), .B0(n2602), .B1(n2601), .Y(n2613) );
  OAI21X1 U1048 ( .A0(n2596), .A1(n2597), .B0(n2604), .Y(n2602) );
  NOR2X1 U1049 ( .A(n2903), .B(n2899), .Y(n2884) );
  OAI21X1 U1050 ( .A0(n1275), .A1(n1278), .B0(n1274), .Y(n1279) );
  OAI21X1 U1051 ( .A0(n2470), .A1(n1270), .B0(n1269), .Y(n1275) );
  AOI2BB1X4 U1052 ( .A0N(n1428), .A1N(n2118), .B0(n2928), .Y(n864) );
  AOI211X1 U1053 ( .A0(n2931), .A1(n257), .B0(n251), .C0(n2928), .Y(n2971) );
  OAI21X1 U1054 ( .A0(n2121), .A1(n1378), .B0(n1433), .Y(n2928) );
  OAI22X1 U1055 ( .A0(n2206), .A1(n2205), .B0(n2204), .B1(n2203), .Y(n2212) );
  NOR3X1 U1056 ( .A(n2647), .B(n2958), .C(n2960), .Y(n2110) );
  AOI21X1 U1057 ( .A0(n1204), .A1(n1206), .B0(n1211), .Y(n1210) );
  NOR3X1 U1058 ( .A(n1206), .B(n1195), .C(n1204), .Y(n1211) );
  NOR3X1 U1059 ( .A(n1632), .B(n1631), .C(n1630), .Y(n1634) );
  NOR2BX1 U1060 ( .AN(n1653), .B(n1665), .Y(n1630) );
  NOR2X1 U1061 ( .A(n2187), .B(n2195), .Y(n2190) );
  NOR3X1 U1062 ( .A(n2179), .B(n76), .C(n2196), .Y(n2187) );
  AOI211X1 U1063 ( .A0(n149), .A1(n277), .B0(n814), .C0(n816), .Y(n783) );
  NAND2X1 U1064 ( .A(global_cntr[17]), .B(n275), .Y(n277) );
  OAI21X1 U1065 ( .A0(N2283), .A1(n41), .B0(n2302), .Y(n2293) );
  NOR2X1 U1066 ( .A(n32), .B(state[2]), .Y(n827) );
  NAND2X1 U1067 ( .A(state[2]), .B(n32), .Y(n833) );
  NOR2X1 U1068 ( .A(state[2]), .B(n185), .Y(n281) );
  NAND2XL U1069 ( .A(n209), .B(\C169/Z_2 ), .Y(n108) );
  NAND2XL U1070 ( .A(\DP_OP_725J1_134_142/I4 ), .B(N744), .Y(n109) );
  OR3X4 U1071 ( .A(n772), .B(n619), .C(n1868), .Y(n209) );
  NOR2X6 U1072 ( .A(read_cntr[0]), .B(n506), .Y(\DP_OP_725J1_134_142/I3 ) );
  NOR4X1 U1073 ( .A(n800), .B(n801), .C(n799), .D(n786), .Y(n819) );
  AOI211X1 U1074 ( .A0(n145), .A1(n262), .B0(n261), .C0(n816), .Y(n799) );
  NAND2X1 U1075 ( .A(write_cntr[9]), .B(n170), .Y(n1883) );
  NOR2X1 U1076 ( .A(n170), .B(write_cntr[9]), .Y(n1884) );
  NAND2X1 U1077 ( .A(n1876), .B(n170), .Y(n1877) );
  AND2X2 U1078 ( .A(n1879), .B(write_cntr[14]), .Y(n170) );
  CLKINVX1 U1079 ( .A(next_cr_x[5]), .Y(n1301) );
  NAND2X2 U1080 ( .A(n1059), .B(n1058), .Y(next_cr_x[5]) );
  CLKINVX1 U1081 ( .A(n765), .Y(sftr_n[1]) );
  AOI31X1 U1082 ( .A0(n765), .A1(n2966), .A2(n2965), .B0(n2964), .Y(n2970) );
  AND2X2 U1083 ( .A(n778), .B(n357), .Y(n765) );
  CLKINVX1 U1084 ( .A(n1071), .Y(n479) );
  NAND2BX1 U1085 ( .AN(n1609), .B(n1611), .Y(n1641) );
  NAND2X1 U1086 ( .A(n1584), .B(n1583), .Y(n1611) );
  OAI21X1 U1087 ( .A0(n1972), .A1(n1971), .B0(n1991), .Y(n1989) );
  NAND2X1 U1088 ( .A(n1971), .B(n1970), .Y(n1991) );
  OAI2BB2X1 U1089 ( .B0(curr_time[12]), .B1(m_1[3]), .A0N(curr_time[12]), 
        .A1N(m_1[3]), .Y(n1022) );
  NAND2X1 U1090 ( .A(n299), .B(n306), .Y(m_1[3]) );
  NAND2X1 U1091 ( .A(n443), .B(n374), .Y(n461) );
  NAND2X1 U1092 ( .A(n373), .B(n375), .Y(n443) );
  AOI22X1 U1093 ( .A0(n1353), .A1(n1352), .B0(n1351), .B1(n1350), .Y(n1354) );
  CLKINVX1 U1094 ( .A(n1348), .Y(n1350) );
  NAND2X1 U1095 ( .A(n1076), .B(write_addr[18]), .Y(n1083) );
  NOR2X1 U1096 ( .A(n1077), .B(n154), .Y(n1076) );
  NAND2X1 U1097 ( .A(n2007), .B(n2006), .Y(n2018) );
  NAND2BX1 U1098 ( .AN(n2198), .B(n2202), .Y(n2225) );
  NAND2X1 U1099 ( .A(n2192), .B(n2191), .Y(n2202) );
  NOR2X1 U1100 ( .A(n2192), .B(n2191), .Y(n2198) );
  NOR3BX1 U1101 ( .AN(n2047), .B(n2056), .C(n2040), .Y(n2048) );
  NOR2X1 U1102 ( .A(n2041), .B(n2040), .Y(n2043) );
  NAND2BX1 U1103 ( .AN(n2033), .B(n2037), .Y(n2040) );
  BUFX4 U1104 ( .A(n614), .Y(n252) );
  NOR2X1 U1105 ( .A(next_work_cntr[1]), .B(n2875), .Y(n2898) );
  OAI2BB2X2 U1106 ( .B0(next_work_cntr[1]), .B1(n2875), .A0N(next_work_cntr[1]), .A1N(n2875), .Y(n2916) );
  NOR2X1 U1107 ( .A(n2893), .B(n2892), .Y(n2875) );
  OAI21X1 U1108 ( .A0(n875), .A1(n874), .B0(n873), .Y(n877) );
  NOR2X1 U1109 ( .A(n867), .B(n175), .Y(n875) );
  NOR2X1 U1110 ( .A(n2088), .B(n2090), .Y(n2089) );
  NOR2X1 U1111 ( .A(n2566), .B(n2567), .Y(n2577) );
  NOR2X1 U1112 ( .A(n2549), .B(n2550), .Y(n2562) );
  OAI221X4 U1113 ( .A0(n2635), .A1(n2634), .B0(n2633), .B1(n2632), .C0(n2631), 
        .Y(n2639) );
  NOR2BX1 U1114 ( .AN(n2625), .B(n2623), .Y(n2632) );
  NOR2X1 U1115 ( .A(n2941), .B(n237), .Y(n2943) );
  NOR2X1 U1116 ( .A(curr_time[9]), .B(n432), .Y(n431) );
  AOI21X1 U1117 ( .A0(n441), .A1(n440), .B0(n390), .Y(n432) );
  NOR2X1 U1118 ( .A(n2531), .B(n2530), .Y(n2542) );
  NAND2X1 U1119 ( .A(n2658), .B(n2708), .Y(n2679) );
  OAI31X1 U1120 ( .A0(n2708), .A1(n2707), .A2(n2706), .B0(n2705), .Y(n2725) );
  NOR2X1 U1121 ( .A(next_work_cntr[9]), .B(n2685), .Y(n2708) );
  NOR2X1 U1122 ( .A(n202), .B(n1878), .Y(n1891) );
  NAND2X1 U1123 ( .A(n2937), .B(cr_read_cntr[5]), .Y(n2939) );
  NOR2X1 U1124 ( .A(n2936), .B(n241), .Y(n2937) );
  AOI2BB2X2 U1125 ( .B0(n2804), .B1(n2803), .A0N(n2804), .A1N(n2803), .Y(n2860) );
  NOR2X1 U1126 ( .A(n2830), .B(n2828), .Y(n2803) );
  NOR2BX1 U1127 ( .AN(n2019), .B(n2020), .Y(n2021) );
  NOR2X1 U1128 ( .A(n2008), .B(n2009), .Y(n2020) );
  NOR2X1 U1129 ( .A(n1874), .B(n1954), .Y(N2900) );
  NOR2BX1 U1130 ( .AN(n1687), .B(N205), .Y(n1682) );
  NAND2BX1 U1131 ( .AN(n1674), .B(n1671), .Y(n1687) );
  OAI21X1 U1132 ( .A0(curr_time[15]), .A1(n804), .B0(n1016), .Y(n1018) );
  OAI21X1 U1133 ( .A0(curr_time[7]), .A1(n805), .B0(n1023), .Y(n1025) );
  OAI21X1 U1134 ( .A0(curr_time[23]), .A1(n803), .B0(n1008), .Y(n1010) );
  NOR2X1 U1135 ( .A(n1699), .B(n1704), .Y(n1708) );
  NOR2X1 U1136 ( .A(n1722), .B(n2965), .Y(n1704) );
  NOR2BX1 U1137 ( .AN(n1174), .B(n1183), .Y(n1180) );
  NOR2X1 U1138 ( .A(n1173), .B(n1172), .Y(n1183) );
  OAI2BB2X2 U1139 ( .B0(n2239), .B1(n2238), .A0N(n2239), .A1N(n2238), .Y(n2259) );
  NOR2X1 U1140 ( .A(n2239), .B(n2238), .Y(n2246) );
  OAI2BB2X1 U1141 ( .B0(n2233), .B1(n2232), .A0N(n2233), .A1N(n2231), .Y(n2238) );
  OAI22X1 U1142 ( .A0(n1235), .A1(n1234), .B0(n1233), .B1(n1232), .Y(n1239) );
  OAI2BB2X1 U1143 ( .B0(n1224), .B1(n1223), .A0N(n1224), .A1N(n1229), .Y(n1234) );
  OAI21X1 U1144 ( .A0(n2770), .A1(n2769), .B0(n2768), .Y(n2791) );
  OAI31X1 U1145 ( .A0(next_work_cntr[6]), .A1(n2741), .A2(n2740), .B0(n2769), 
        .Y(n2768) );
  OAI21X1 U1146 ( .A0(n2742), .A1(n2739), .B0(n2738), .Y(n2769) );
  OAI21X1 U1147 ( .A0(n2719), .A1(n2718), .B0(n2717), .Y(n2742) );
  NAND2X1 U1148 ( .A(n2213), .B(n2212), .Y(n2224) );
  NOR2X1 U1149 ( .A(n2213), .B(n2212), .Y(n2222) );
  OAI21X1 U1150 ( .A0(n2194), .A1(n2670), .B0(n2193), .Y(n2213) );
  OAI22X1 U1151 ( .A0(n1128), .A1(n1127), .B0(n1129), .B1(n1126), .Y(n1143) );
  NAND2X2 U1152 ( .A(n1130), .B(n1129), .Y(\intadd_3/A[0] ) );
  OAI21X1 U1153 ( .A0(n1117), .A1(n1116), .B0(n1115), .Y(n1129) );
  OAI21X1 U1154 ( .A0(n2353), .A1(n2352), .B0(n2351), .Y(n2359) );
  OAI21X1 U1155 ( .A0(n2410), .A1(n2409), .B0(n2408), .Y(n2416) );
  OAI21X1 U1156 ( .A0(n2671), .A1(n2391), .B0(n2390), .Y(n2397) );
  OAI21X1 U1157 ( .A0(n2430), .A1(n2429), .B0(n2428), .Y(n2436) );
  OAI2BB2X1 U1158 ( .B0(n1388), .B1(n88), .A0N(n1388), .A1N(n88), .Y(n1386) );
  NAND2X1 U1159 ( .A(n1074), .B(n89), .Y(n1388) );
  OAI21X1 U1160 ( .A0(n1573), .A1(n61), .B0(n1571), .Y(n1615) );
  OAI21X1 U1161 ( .A0(n1440), .A1(n188), .B0(n1442), .Y(n1459) );
  OAI2BB2X1 U1162 ( .B0(n1073), .B1(n102), .A0N(n1073), .A1N(n102), .Y(n1377)
         );
  OAI21X1 U1163 ( .A0(n1848), .A1(n1847), .B0(n1846), .Y(n1850) );
  OAI22X1 U1164 ( .A0(n1882), .A1(n1881), .B0(n1889), .B1(n1888), .Y(n1902) );
  OAI22X1 U1165 ( .A0(n1064), .A1(n1063), .B0(cr_read_cntr[6]), .B1(n1062), 
        .Y(n1065) );
  OAI22X1 U1166 ( .A0(n1670), .A1(n1669), .B0(n1668), .B1(n1667), .Y(n1676) );
  AOI2BB2X2 U1167 ( .B0(n1020), .B1(n387), .A0N(n386), .A1N(n1021), .Y(n442)
         );
  NOR3X1 U1168 ( .A(n1259), .B(n1255), .C(n1258), .Y(n1264) );
  OAI22X1 U1169 ( .A0(n1252), .A1(n1250), .B0(n1249), .B1(n1248), .Y(n1258) );
  AOI211X1 U1170 ( .A0(n139), .A1(n818), .B0(n265), .C0(n266), .Y(n792) );
  NOR3BX1 U1171 ( .AN(n1123), .B(n1103), .C(n2139), .Y(n1109) );
  OAI22X1 U1172 ( .A0(n2135), .A1(n1301), .B0(n1057), .B1(next_cr_x[5]), .Y(
        n1103) );
  CLKINVX1 U1173 ( .A(n2142), .Y(n881) );
  OAI2BB2X1 U1174 ( .B0(n2688), .B1(n2687), .A0N(n2688), .A1N(n2687), .Y(n2700) );
  OAI31X4 U1175 ( .A0(n2661), .A1(n2660), .A2(n2662), .B0(n2659), .Y(n2687) );
  OAI31X1 U1176 ( .A0(n83), .A1(n969), .A2(n968), .B0(n967), .Y(n977) );
  OAI2BB2X1 U1177 ( .B0(n1012), .B1(n1011), .A0N(n1012), .A1N(n1011), .Y(n1013) );
  XOR2X1 U1178 ( .A(n46), .B(curr_time[20]), .Y(n1011) );
  OAI2BB2X2 U1179 ( .B0(n1027), .B1(n1026), .A0N(n1027), .A1N(n1026), .Y(n1028) );
  XNOR2X1 U1180 ( .A(\h_1[2] ), .B(n297), .Y(n1014) );
  NAND2X1 U1181 ( .A(n405), .B(n404), .Y(\h_1[2] ) );
  XOR2X1 U1182 ( .A(\s_1[2] ), .B(curr_time[3]), .Y(n1030) );
  NOR2X1 U1183 ( .A(n2860), .B(n2878), .Y(n2864) );
  OAI31X1 U1184 ( .A0(n1348), .A1(n1351), .A2(n1349), .B0(n1347), .Y(n1356) );
  NOR2X2 U1185 ( .A(n944), .B(n943), .Y(n1348) );
  CLKINVX1 U1186 ( .A(n2686), .Y(next_work_cntr[9]) );
  NAND2X1 U1187 ( .A(n2151), .B(n2686), .Y(n2218) );
  OA21X1 U1188 ( .A0(n2151), .A1(n2686), .B0(n2218), .Y(n2239) );
  OAI2BB2X2 U1189 ( .B0(n2686), .B1(n2685), .A0N(n2686), .A1N(n2685), .Y(n2731) );
  CLKINVX1 U1190 ( .A(n1283), .Y(n1415) );
  NAND2X1 U1191 ( .A(n1154), .B(n1153), .Y(n1283) );
  NOR2X2 U1192 ( .A(n41), .B(n2372), .Y(next_work_cntr[13]) );
  OAI21X1 U1193 ( .A0(n2372), .A1(n2371), .B0(n2370), .Y(n2378) );
  CLKINVX1 U1194 ( .A(n2652), .Y(n2372) );
  AND2X2 U1195 ( .A(n1918), .B(n2131), .Y(n1930) );
  CLKINVX1 U1196 ( .A(n2131), .Y(n806) );
  NOR2X2 U1197 ( .A(n2131), .B(n465), .Y(n470) );
  NAND2X1 U1198 ( .A(n257), .B(n2333), .Y(n2664) );
  CLKINVX1 U1199 ( .A(n2312), .Y(n2333) );
  CLKINVX1 U1200 ( .A(n778), .Y(n1721) );
  NOR2X2 U1201 ( .A(state[0]), .B(n282), .Y(n778) );
  NOR3X1 U1202 ( .A(n2951), .B(n2950), .C(n2949), .Y(n2952) );
  NAND2X1 U1203 ( .A(n796), .B(n2321), .Y(n2949) );
  NOR2X2 U1204 ( .A(n169), .B(n233), .Y(n1713) );
  NOR2X2 U1205 ( .A(n2649), .B(n2653), .Y(n2678) );
  NAND2X1 U1206 ( .A(next_work_cntr[19]), .B(n2655), .Y(n2653) );
  OAI2BB2X2 U1207 ( .B0(n1569), .B1(n1568), .A0N(n1569), .A1N(n1568), .Y(n1605) );
  NOR2BX2 U1208 ( .AN(n1548), .B(n1549), .Y(n1569) );
  NOR2X2 U1209 ( .A(n1706), .B(n207), .Y(n771) );
  CLKINVX1 U1210 ( .A(n1684), .Y(n1706) );
  NAND2X2 U1211 ( .A(n1721), .B(n771), .Y(n1868) );
  NAND2BX1 U1212 ( .AN(n2276), .B(n2272), .Y(n2279) );
  NOR2X2 U1213 ( .A(n2265), .B(n2264), .Y(n2276) );
  NOR2BX2 U1214 ( .AN(n1598), .B(n1599), .Y(n1629) );
  NAND2X1 U1215 ( .A(n164), .B(n1570), .Y(n1598) );
  NOR2X1 U1216 ( .A(n164), .B(n1570), .Y(n1599) );
  NOR2XL U1217 ( .A(n2034), .B(n2014), .Y(n111) );
  NOR2XL U1218 ( .A(work_cntr[9]), .B(n2014), .Y(n112) );
  NOR2X4 U1219 ( .A(work_cntr[9]), .B(n2034), .Y(n2014) );
  NAND2BX1 U1220 ( .AN(n110), .B(n2036), .Y(n2041) );
  NAND2X1 U1221 ( .A(n2035), .B(n193), .Y(n2034) );
  NOR2X2 U1222 ( .A(n842), .B(n849), .Y(n848) );
  NAND2X1 U1223 ( .A(write_cntr[10]), .B(n851), .Y(n849) );
  NOR2BX2 U1224 ( .AN(n2055), .B(n2050), .Y(n2061) );
  OAI21X1 U1225 ( .A0(n2048), .A1(n2046), .B0(n2047), .Y(n2055) );
  BUFX2 U1226 ( .A(n2023), .Y(n113) );
  AOI22X1 U1227 ( .A0(n2025), .A1(n2024), .B0(n113), .B1(n2022), .Y(n2027) );
  NAND2X1 U1228 ( .A(n114), .B(n115), .Y(n1913) );
  CLKINVX1 U1229 ( .A(n1894), .Y(n116) );
  INVXL U1230 ( .A(n1895), .Y(n117) );
  NAND2XL U1231 ( .A(n1895), .B(n1894), .Y(n114) );
  NAND2X1 U1232 ( .A(n116), .B(n117), .Y(n115) );
  OAI2BB2X1 U1233 ( .B0(n1913), .B1(n1912), .A0N(n1913), .A1N(n1912), .Y(n1921) );
  NOR2BX2 U1234 ( .AN(n1883), .B(n1884), .Y(n1895) );
  NOR2X1 U1235 ( .A(n2098), .B(n2969), .Y(expand_sel[1]) );
  NOR2BX2 U1236 ( .AN(n1908), .B(n1909), .Y(n1926) );
  NOR2X1 U1237 ( .A(write_cntr[7]), .B(n1950), .Y(n1909) );
  NAND2X1 U1238 ( .A(write_cntr[7]), .B(n1950), .Y(n1908) );
  NOR2BX2 U1239 ( .AN(n2241), .B(n2237), .Y(n2247) );
  NOR2X1 U1240 ( .A(n2229), .B(n2228), .Y(n2237) );
  NAND2X1 U1241 ( .A(n2229), .B(n2228), .Y(n2241) );
  AOI22X2 U1242 ( .A0(n2927), .A1(n2926), .B0(n777), .B1(n2925), .Y(n2931) );
  NAND2X1 U1243 ( .A(n118), .B(n119), .Y(n1650) );
  CLKINVX1 U1244 ( .A(n1581), .Y(n120) );
  INVXL U1245 ( .A(n1580), .Y(n121) );
  NAND2XL U1246 ( .A(n1580), .B(n1581), .Y(n118) );
  NAND2X1 U1247 ( .A(n120), .B(n121), .Y(n119) );
  NOR2X1 U1248 ( .A(n1574), .B(n1598), .Y(n1581) );
  OAI2BB2X2 U1249 ( .B0(n1551), .B1(n1550), .A0N(n1551), .A1N(n1550), .Y(n1580) );
  NAND2X1 U1250 ( .A(n2792), .B(n2791), .Y(n2787) );
  CLKINVX1 U1251 ( .A(n2771), .Y(next_work_cntr[5]) );
  OAI21X1 U1252 ( .A0(n1015), .A1(n410), .B0(n415), .Y(n419) );
  NAND2X1 U1253 ( .A(n122), .B(n123), .Y(n1898) );
  CLKINVX1 U1254 ( .A(n1885), .Y(n124) );
  NAND2XL U1255 ( .A(write_cntr[10]), .B(n1885), .Y(n122) );
  NAND2X1 U1256 ( .A(n124), .B(n204), .Y(n123) );
  NAND2X1 U1257 ( .A(n125), .B(n126), .Y(n1931) );
  CLKINVX1 U1258 ( .A(n1910), .Y(n127) );
  INVXL U1259 ( .A(n1911), .Y(n128) );
  NAND2XL U1260 ( .A(n1911), .B(n1910), .Y(n125) );
  NAND2X1 U1261 ( .A(n127), .B(n128), .Y(n126) );
  OAI21X1 U1262 ( .A0(n1909), .A1(n1924), .B0(n1908), .Y(n1910) );
  NOR2BX2 U1263 ( .AN(n1892), .B(n1893), .Y(n1911) );
  NOR2X1 U1264 ( .A(n1557), .B(n1578), .Y(n1559) );
  NOR2X1 U1265 ( .A(n1557), .B(n1497), .Y(n1519) );
  NOR2X1 U1266 ( .A(n1557), .B(n1554), .Y(n1534) );
  AOI2BB2X2 U1267 ( .B0(n180), .B1(n1482), .A0N(n180), .A1N(n1482), .Y(n1557)
         );
  CLKINVX1 U1268 ( .A(n2493), .Y(n2486) );
  NOR2X2 U1269 ( .A(n2099), .B(n2120), .Y(n2493) );
  CLKINVX1 U1270 ( .A(n1335), .Y(n1334) );
  NOR2X2 U1271 ( .A(n905), .B(n908), .Y(n1335) );
  CLKINVX1 U1272 ( .A(n1444), .Y(n1960) );
  OA21X1 U1273 ( .A0(n2154), .A1(n2153), .B0(n2167), .Y(n2179) );
  NOR2X2 U1274 ( .A(n2656), .B(n2167), .Y(n2157) );
  NAND2X2 U1275 ( .A(n2154), .B(n2153), .Y(n2167) );
  AND2X2 U1276 ( .A(n1002), .B(n996), .Y(n1310) );
  NAND2X1 U1277 ( .A(work_cntr[17]), .B(n1032), .Y(n1031) );
  OAI21X1 U1278 ( .A0(work_cntr[17]), .A1(n1032), .B0(n1031), .Y(n2312) );
  CLKINVX1 U1279 ( .A(n2751), .Y(next_work_cntr[6]) );
  NOR2X2 U1280 ( .A(n985), .B(n990), .Y(n1319) );
  NOR2X2 U1281 ( .A(n2851), .B(n2849), .Y(n2882) );
  NOR2X1 U1282 ( .A(n768), .B(n364), .Y(n467) );
  NOR2X2 U1283 ( .A(n2130), .B(n356), .Y(n768) );
  NAND2X1 U1284 ( .A(n1683), .B(write_addr[8]), .Y(n1366) );
  CLKAND2X3 U1285 ( .A(\next_write_addr_w[0] ), .B(n1683), .Y(n772) );
  NOR2BX2 U1286 ( .AN(n1079), .B(n168), .Y(n1683) );
  OAI2BB2X2 U1287 ( .B0(n2684), .B1(n2683), .A0N(n2684), .A1N(n2683), .Y(n2727) );
  NOR2BX1 U1288 ( .AN(n2679), .B(n2678), .Y(n2683) );
  NOR2BX2 U1289 ( .AN(n1516), .B(n1515), .Y(n1512) );
  OAI21X1 U1290 ( .A0(n2801), .A1(n2800), .B0(n2799), .Y(n2821) );
  NOR2X1 U1291 ( .A(n2813), .B(n2800), .Y(n2788) );
  NOR2X1 U1292 ( .A(n2800), .B(n2801), .Y(n2773) );
  OAI2BB2X2 U1293 ( .B0(n2749), .B1(n2748), .A0N(n2749), .A1N(n2748), .Y(n2800) );
  OAI31X4 U1294 ( .A0(n2797), .A1(n2811), .A2(n2810), .B0(n2796), .Y(n2838) );
  NAND2X1 U1295 ( .A(n2811), .B(n2810), .Y(n2835) );
  OAI2BB2X2 U1296 ( .B0(n2782), .B1(n80), .A0N(n2782), .A1N(n80), .Y(n2811) );
  NAND2X1 U1297 ( .A(n2755), .B(n2754), .Y(n2782) );
  NAND2X1 U1298 ( .A(n2760), .B(n2761), .Y(n2777) );
  OAI31X4 U1299 ( .A0(n2762), .A1(n2761), .A2(n2760), .B0(n2759), .Y(n2813) );
  OAI2BB2X2 U1300 ( .B0(n2712), .B1(n2711), .A0N(n2712), .A1N(n2711), .Y(n2761) );
  NOR2X1 U1301 ( .A(n2710), .B(n2709), .Y(n2711) );
  NOR2X2 U1302 ( .A(n366), .B(n365), .Y(n469) );
  NOR2X1 U1303 ( .A(n1587), .B(n1586), .Y(n1558) );
  NOR2X1 U1304 ( .A(n1587), .B(n1585), .Y(n1584) );
  OAI2BB2X2 U1305 ( .B0(n82), .B1(n1528), .A0N(n82), .A1N(n1528), .Y(n1587) );
  NAND2X1 U1306 ( .A(n1526), .B(n1525), .Y(n1528) );
  NOR2X2 U1307 ( .A(n41), .B(n2394), .Y(next_work_cntr[10]) );
  OA21X1 U1308 ( .A0(n2394), .A1(n2400), .B0(n2395), .Y(n2404) );
  CLKINVX1 U1309 ( .A(n2394), .Y(n2649) );
  OAI21X2 U1310 ( .A0(work_cntr[10]), .A1(n1040), .B0(n1039), .Y(n2394) );
  NAND2X1 U1311 ( .A(work_cntr[10]), .B(n1040), .Y(n1039) );
  NOR2X1 U1312 ( .A(n187), .B(n1041), .Y(n1040) );
  OAI21X2 U1313 ( .A0(n63), .A1(write_addr[16]), .B0(n1077), .Y(n1396) );
  NOR3BX1 U1314 ( .AN(n1397), .B(n154), .C(n1396), .Y(n1405) );
  OAI21X1 U1315 ( .A0(n2336), .A1(n2344), .B0(n2340), .Y(n2342) );
  OAI21X2 U1316 ( .A0(work_cntr[16]), .A1(n1034), .B0(n1033), .Y(n2336) );
  OAI22X2 U1317 ( .A0(n2654), .A1(n2308), .B0(next_work_cntr[19]), .B1(n2155), 
        .Y(n2163) );
  CLKINVX1 U1318 ( .A(n1133), .Y(n2134) );
  AOI21X2 U1319 ( .A0(n166), .A1(n952), .B0(n951), .Y(n1133) );
  NAND2X2 U1320 ( .A(n777), .B(n1406), .Y(n1398) );
  CLKINVX1 U1321 ( .A(n1404), .Y(n1406) );
  AND2X2 U1322 ( .A(n257), .B(n283), .Y(n777) );
  CLKINVX1 U1323 ( .A(n1322), .Y(n1325) );
  NOR2X2 U1324 ( .A(n876), .B(n877), .Y(n1322) );
  OAI2BB2X1 U1325 ( .B0(work_cntr[11]), .B1(n2541), .A0N(work_cntr[11]), .A1N(
        n2541), .Y(n2016) );
  OAI31X4 U1326 ( .A0(n2765), .A1(n2764), .A2(n2774), .B0(n2763), .Y(n2822) );
  NAND2X1 U1327 ( .A(n2751), .B(n2750), .Y(n2774) );
  NOR2X2 U1328 ( .A(n41), .B(n2482), .Y(next_work_cntr[2]) );
  NOR2X2 U1329 ( .A(work_cntr[4]), .B(work_cntr[5]), .Y(n2500) );
  OAI2BB2X1 U1330 ( .B0(n1521), .B1(n1520), .A0N(n1562), .A1N(n1563), .Y(n1522) );
  NOR3BX1 U1331 ( .AN(n1485), .B(n1521), .C(n1496), .Y(n1509) );
  NOR2X1 U1332 ( .A(n256), .B(n1521), .Y(n1465) );
  NOR2X1 U1333 ( .A(n1521), .B(n1500), .Y(n1486) );
  OAI2BB2X2 U1334 ( .B0(n1521), .B1(n1502), .A0N(n1521), .A1N(n1502), .Y(n1562) );
  OAI21X2 U1335 ( .A0(n1441), .A1(n184), .B0(n1471), .Y(n1521) );
  NAND2X1 U1336 ( .A(n1441), .B(n184), .Y(n1471) );
  OAI21X1 U1337 ( .A0(n1346), .A1(n1345), .B0(n1344), .Y(n1349) );
  CLKINVX2 U1338 ( .A(n712), .Y(n707) );
  NAND2X2 U1339 ( .A(read_cntr[0]), .B(n1867), .Y(n712) );
  AND2X2 U1340 ( .A(n1475), .B(n2502), .Y(n1460) );
  OA21X2 U1341 ( .A0(n2502), .A1(n1747), .B0(n1742), .Y(n1750) );
  OAI21X2 U1342 ( .A0(n1187), .A1(n2502), .B0(n1186), .Y(n1200) );
  INVX3 U1343 ( .A(n256), .Y(n2502) );
  CLKINVX1 U1344 ( .A(n1308), .Y(n1298) );
  NAND2X2 U1345 ( .A(n1098), .B(n1097), .Y(n1308) );
  CLKBUFX3 U1346 ( .A(work_cntr[7]), .Y(n129) );
  OAI21X2 U1347 ( .A0(n129), .A1(n1044), .B0(n1043), .Y(n2430) );
  NOR2X1 U1348 ( .A(n129), .B(n1226), .Y(n1227) );
  AOI21X2 U1349 ( .A0(n129), .A1(n1958), .B0(n2035), .Y(n2051) );
  NOR2X1 U1350 ( .A(n129), .B(n1958), .Y(n2035) );
  AOI2BB2X2 U1351 ( .B0(n129), .B1(n1512), .A0N(n129), .A1N(n1512), .Y(n1551)
         );
  NOR2X1 U1352 ( .A(n129), .B(n1512), .Y(n1527) );
  CLKINVX2 U1353 ( .A(n861), .Y(next_cr_x[6]) );
  CLKINVX1 U1354 ( .A(n703), .Y(n701) );
  OR2X4 U1355 ( .A(n623), .B(n710), .Y(n703) );
  NOR2BX1 U1356 ( .AN(n950), .B(n1135), .Y(n948) );
  CLKINVX1 U1357 ( .A(n1135), .Y(n2138) );
  OAI32X4 U1358 ( .A0(write_cntr[5]), .A1(n166), .A2(n952), .B0(n951), .B1(
        n198), .Y(n1135) );
  BUFX2 U1359 ( .A(n1340), .Y(n130) );
  NOR2X1 U1360 ( .A(n924), .B(n130), .Y(n923) );
  OAI2BB2X1 U1361 ( .B0(n1341), .B1(n130), .A0N(n1341), .A1N(n1339), .Y(n1346)
         );
  NOR2X1 U1362 ( .A(n2930), .B(n1428), .Y(n132) );
  CLKINVX1 U1363 ( .A(n2929), .Y(n133) );
  AOI32X4 U1364 ( .A0(n204), .A1(n131), .A2(n851), .B0(n852), .B1(
        write_cntr[10]), .Y(n2142) );
  AOI32X4 U1365 ( .A0(n907), .A1(n196), .A2(n131), .B0(write_cntr[7]), .B1(
        n906), .Y(n2140) );
  AOI21X1 U1366 ( .A0(n131), .A1(n932), .B0(n975), .Y(n951) );
  CLKINVX1 U1367 ( .A(n251), .Y(n1428) );
  NAND2X2 U1368 ( .A(n1962), .B(n152), .Y(n2955) );
  INVX3 U1369 ( .A(n1434), .Y(n1431) );
  BUFX16 U1370 ( .A(n2976), .Y(cr_a[4]) );
  NOR2BX1 U1371 ( .AN(N1457), .B(n2969), .Y(n2976) );
  OR2X4 U1372 ( .A(n721), .B(n720), .Y(n759) );
  INVX3 U1373 ( .A(n769), .Y(n597) );
  AND2X2 U1374 ( .A(n1695), .B(n771), .Y(n769) );
  CLKINVX1 U1375 ( .A(n612), .Y(n615) );
  CLKAND2X3 U1376 ( .A(n512), .B(n511), .Y(n612) );
  AND2X2 U1377 ( .A(n2126), .B(n322), .Y(n2972) );
  INVX16 U1378 ( .A(n2972), .Y(im_wen_n) );
  INVX4 U1379 ( .A(n780), .Y(n717) );
  NOR2X6 U1380 ( .A(n718), .B(n622), .Y(\DP_OP_725J1_134_142/I7 ) );
  AOI22XL U1381 ( .A0(n209), .A1(\C169/Z_0 ), .B0(\DP_OP_725J1_134_142/I4 ), 
        .B1(N742), .Y(\DP_OP_725J1_134_142/n144 ) );
  AOI22XL U1382 ( .A0(n209), .A1(\C169/Z_1 ), .B0(\DP_OP_725J1_134_142/I4 ), 
        .B1(N743), .Y(\DP_OP_725J1_134_142/n142 ) );
  AOI22XL U1383 ( .A0(n209), .A1(\C169/Z_3 ), .B0(\DP_OP_725J1_134_142/I4 ), 
        .B1(N745), .Y(\DP_OP_725J1_134_142/n136 ) );
  AOI22XL U1384 ( .A0(n209), .A1(\C169/Z_4 ), .B0(\DP_OP_725J1_134_142/I4 ), 
        .B1(N746), .Y(\DP_OP_725J1_134_142/n133 ) );
  AOI22XL U1385 ( .A0(n209), .A1(\C169/Z_5 ), .B0(\DP_OP_725J1_134_142/I4 ), 
        .B1(N747), .Y(\DP_OP_725J1_134_142/n130 ) );
  NOR2X6 U1386 ( .A(n171), .B(n506), .Y(\DP_OP_725J1_134_142/I4 ) );
  NOR3X6 U1387 ( .A(n772), .B(n1868), .C(n1869), .Y(\DP_OP_725J1_134_142/I2 )
         );
  AOI22XL U1388 ( .A0(n173), .A1(\DP_OP_725J1_134_142/I3 ), .B0(n173), .B1(
        \DP_OP_725J1_134_142/I2 ), .Y(\DP_OP_725J1_134_142/n143 ) );
  NAND2XL U1389 ( .A(N622), .B(\DP_OP_725J1_134_142/I2 ), .Y(
        \DP_OP_725J1_134_142/n141 ) );
  NAND2XL U1390 ( .A(N623), .B(\DP_OP_725J1_134_142/I2 ), .Y(
        \DP_OP_725J1_134_142/n138 ) );
  NAND2XL U1391 ( .A(N624), .B(\DP_OP_725J1_134_142/I2 ), .Y(
        \DP_OP_725J1_134_142/n135 ) );
  NAND2XL U1392 ( .A(N625), .B(\DP_OP_725J1_134_142/I2 ), .Y(
        \DP_OP_725J1_134_142/n132 ) );
  NAND2XL U1393 ( .A(N626), .B(\DP_OP_725J1_134_142/I2 ), .Y(
        \DP_OP_725J1_134_142/n129 ) );
  NAND2X1 U1394 ( .A(global_cntr[2]), .B(n1873), .Y(n1954) );
  INVXL U1395 ( .A(n798), .Y(n1953) );
  NOR2X2 U1396 ( .A(n1874), .B(n1952), .Y(N2858) );
  NAND3X2 U1397 ( .A(n32), .B(n163), .C(n190), .Y(N2902) );
  INVXL U1398 ( .A(n2820), .Y(next_work_cntr[3]) );
  INVXL U1399 ( .A(n2670), .Y(next_work_cntr[12]) );
  NAND2XL U1400 ( .A(curr_photo[0]), .B(n243), .Y(n360) );
  NOR2XL U1401 ( .A(curr_photo[0]), .B(n2953), .Y(n2951) );
  NOR2XL U1402 ( .A(n2949), .B(n2950), .Y(n2946) );
  NOR2BXL U1403 ( .AN(N1456), .B(n2969), .Y(n2977) );
  NOR2BXL U1404 ( .AN(N1458), .B(n2969), .Y(n2975) );
  NOR2BXL U1405 ( .AN(N1459), .B(n2969), .Y(n2974) );
  NOR2BXL U1406 ( .AN(N1460), .B(n2969), .Y(n2973) );
  OAI211XL U1407 ( .A0(n425), .A1(n419), .B0(n473), .C0(n418), .Y(n420) );
  INVXL U1408 ( .A(n460), .Y(n417) );
  AOI211XL U1409 ( .A0(n469), .A1(n402), .B0(n401), .C0(n400), .Y(n421) );
  AOI211XL U1410 ( .A0(n431), .A1(n399), .B0(n448), .C0(n398), .Y(n400) );
  AOI21XL U1411 ( .A0(n399), .A1(n458), .B0(n431), .Y(n398) );
  XNOR2XL U1412 ( .A(n380), .B(n379), .Y(n383) );
  NAND2XL U1413 ( .A(n461), .B(n429), .Y(n380) );
  INVXL U1414 ( .A(m_1[3]), .Y(n422) );
  NAND3XL U1415 ( .A(n439), .B(n438), .C(n437), .Y(\C1/Z_2 ) );
  AOI22XL U1416 ( .A0(n471), .A1(n436), .B0(n469), .B1(\s_1[2] ), .Y(n437) );
  INVXL U1417 ( .A(n431), .Y(n435) );
  AOI22XL U1418 ( .A0(n470), .A1(\h_1[2] ), .B0(n472), .B1(n430), .Y(n438) );
  NOR2XL U1419 ( .A(curr_time[1]), .B(n443), .Y(n427) );
  AOI22XL U1420 ( .A0(n459), .A1(m_1[2]), .B0(n473), .B1(n426), .Y(n439) );
  NOR2XL U1421 ( .A(curr_time[17]), .B(n452), .Y(n423) );
  INVXL U1422 ( .A(n407), .Y(n406) );
  INVXL U1423 ( .A(n465), .Y(n466) );
  OAI211XL U1424 ( .A0(curr_time[17]), .A1(n454), .B0(n473), .C0(n453), .Y(
        n455) );
  NAND2XL U1425 ( .A(curr_time[17]), .B(n460), .Y(n453) );
  INVXL U1426 ( .A(n452), .Y(n454) );
  AOI211XL U1427 ( .A0(n469), .A1(n451), .B0(n450), .C0(n449), .Y(n456) );
  AOI211XL U1428 ( .A0(curr_time[9]), .A1(n458), .B0(n448), .C0(n447), .Y(n449) );
  NOR2XL U1429 ( .A(curr_time[9]), .B(n446), .Y(n447) );
  MXI2XL U1430 ( .A(n443), .B(n461), .S0(curr_time[1]), .Y(n445) );
  NAND2XL U1431 ( .A(n376), .B(n375), .Y(n451) );
  INVXL U1432 ( .A(n1070), .Y(n478) );
  INVXL U1433 ( .A(n473), .Y(n475) );
  NOR4XL U1434 ( .A(n472), .B(n471), .C(n470), .D(n469), .Y(n476) );
  NAND3XL U1435 ( .A(n464), .B(n463), .C(n462), .Y(\C1/Z_0 ) );
  AOI22XL U1436 ( .A0(\m_0[0] ), .A1(n471), .B0(n469), .B1(n461), .Y(n462) );
  NAND2BXL U1437 ( .AN(n1028), .B(n1029), .Y(n375) );
  OAI211XL U1438 ( .A0(n378), .A1(n372), .B0(n1028), .C0(n376), .Y(n373) );
  INVXL U1439 ( .A(n368), .Y(n370) );
  INVXL U1440 ( .A(n367), .Y(n371) );
  INVXL U1441 ( .A(curr_time[2]), .Y(n372) );
  INVXL U1442 ( .A(n1030), .Y(n378) );
  INVXL U1443 ( .A(n319), .Y(n320) );
  INVXL U1444 ( .A(curr_time[6]), .Y(n317) );
  NAND3XL U1445 ( .A(n316), .B(n315), .C(n314), .Y(n369) );
  NAND2XL U1446 ( .A(n367), .B(n319), .Y(n314) );
  NAND2XL U1447 ( .A(n313), .B(n1025), .Y(n367) );
  NAND2XL U1448 ( .A(n402), .B(n312), .Y(n313) );
  NAND2BXL U1449 ( .AN(n1025), .B(curr_time[4]), .Y(n315) );
  NAND2BXL U1450 ( .AN(n1026), .B(n311), .Y(n316) );
  INVXL U1451 ( .A(curr_time[3]), .Y(n311) );
  NOR2XL U1452 ( .A(curr_time[5]), .B(curr_time[6]), .Y(n1024) );
  NAND3XL U1453 ( .A(n318), .B(curr_time[6]), .C(n309), .Y(n310) );
  NAND2BXL U1454 ( .AN(curr_time[5]), .B(curr_time[7]), .Y(n309) );
  NAND2BXL U1455 ( .AN(n1025), .B(n312), .Y(n318) );
  INVXL U1456 ( .A(curr_time[4]), .Y(n312) );
  NAND3XL U1457 ( .A(curr_time[7]), .B(curr_time[6]), .C(n805), .Y(n1023) );
  INVXL U1458 ( .A(curr_time[5]), .Y(n805) );
  INVXL U1459 ( .A(n467), .Y(n365) );
  INVXL U1460 ( .A(n448), .Y(n471) );
  AOI22XL U1461 ( .A0(n470), .A1(n460), .B0(n472), .B1(\s_0[0] ), .Y(n463) );
  NAND2XL U1462 ( .A(n2131), .B(n381), .Y(n364) );
  OAI211XL U1463 ( .A0(n412), .A1(n411), .B0(n1013), .C0(n410), .Y(n414) );
  INVXL U1464 ( .A(n1014), .Y(n412) );
  NAND2XL U1465 ( .A(n1014), .B(n407), .Y(n415) );
  NAND2XL U1466 ( .A(n444), .B(n411), .Y(n407) );
  INVXL U1467 ( .A(curr_time[18]), .Y(n411) );
  NAND2XL U1468 ( .A(n410), .B(n413), .Y(n444) );
  NAND2BXL U1469 ( .AN(n1013), .B(n1015), .Y(n413) );
  INVXL U1470 ( .A(n294), .Y(n295) );
  NOR2XL U1471 ( .A(n293), .B(n292), .Y(n296) );
  INVXL U1472 ( .A(curr_time[22]), .Y(n292) );
  NAND3XL U1473 ( .A(n291), .B(n290), .C(n289), .Y(n405) );
  NAND2XL U1474 ( .A(n403), .B(n294), .Y(n289) );
  NAND2XL U1475 ( .A(n288), .B(n1010), .Y(n403) );
  NAND2XL U1476 ( .A(n46), .B(n287), .Y(n288) );
  NAND2BXL U1477 ( .AN(n1010), .B(curr_time[20]), .Y(n290) );
  NAND2BXL U1478 ( .AN(n1011), .B(n297), .Y(n291) );
  INVXL U1479 ( .A(curr_time[19]), .Y(n297) );
  NAND2XL U1480 ( .A(curr_time[23]), .B(n1009), .Y(n294) );
  NOR2XL U1481 ( .A(curr_time[21]), .B(curr_time[22]), .Y(n1009) );
  NAND3XL U1482 ( .A(n293), .B(curr_time[22]), .C(n285), .Y(n286) );
  NAND2BXL U1483 ( .AN(curr_time[21]), .B(curr_time[23]), .Y(n285) );
  NAND2BXL U1484 ( .AN(n1010), .B(n287), .Y(n293) );
  INVXL U1485 ( .A(curr_time[20]), .Y(n287) );
  NAND3XL U1486 ( .A(curr_time[23]), .B(curr_time[22]), .C(n803), .Y(n1008) );
  INVXL U1487 ( .A(curr_time[21]), .Y(n803) );
  INVXL U1488 ( .A(curr_time[17]), .Y(n416) );
  AOI22XL U1489 ( .A0(n459), .A1(n458), .B0(\h_0[0] ), .B1(n473), .Y(n464) );
  INVXL U1490 ( .A(curr_time[10]), .Y(n389) );
  NOR2XL U1491 ( .A(n391), .B(curr_time[10]), .Y(n388) );
  NAND3XL U1492 ( .A(n397), .B(n442), .C(n440), .Y(n394) );
  NAND2XL U1493 ( .A(n392), .B(n391), .Y(n395) );
  INVXL U1494 ( .A(n442), .Y(n391) );
  INVXL U1495 ( .A(n397), .Y(n392) );
  INVXL U1496 ( .A(n1022), .Y(n387) );
  NAND2XL U1497 ( .A(n1019), .B(m_1[2]), .Y(n1020) );
  INVXL U1498 ( .A(n306), .Y(n307) );
  NOR2XL U1499 ( .A(n305), .B(n304), .Y(n308) );
  INVXL U1500 ( .A(curr_time[14]), .Y(n304) );
  NAND3XL U1501 ( .A(n303), .B(n1021), .C(n302), .Y(n384) );
  NAND2BXL U1502 ( .AN(n1018), .B(curr_time[12]), .Y(n302) );
  NAND2XL U1503 ( .A(n1022), .B(n1019), .Y(n1021) );
  INVXL U1504 ( .A(curr_time[11]), .Y(n1019) );
  NAND2XL U1505 ( .A(n385), .B(n306), .Y(n303) );
  NAND2XL U1506 ( .A(n301), .B(n1018), .Y(n385) );
  NAND2XL U1507 ( .A(m_1[3]), .B(n300), .Y(n301) );
  NOR2XL U1508 ( .A(curr_time[13]), .B(curr_time[14]), .Y(n1017) );
  NAND3XL U1509 ( .A(n305), .B(curr_time[14]), .C(n298), .Y(n299) );
  NAND2BXL U1510 ( .AN(curr_time[13]), .B(curr_time[15]), .Y(n298) );
  NAND2BXL U1511 ( .AN(n1018), .B(n300), .Y(n305) );
  INVXL U1512 ( .A(curr_time[12]), .Y(n300) );
  NAND3XL U1513 ( .A(curr_time[15]), .B(curr_time[14]), .C(n804), .Y(n1016) );
  INVXL U1514 ( .A(curr_time[13]), .Y(n804) );
  INVXL U1515 ( .A(n474), .Y(n459) );
  INVXL U1516 ( .A(n768), .Y(n408) );
  NAND3XL U1517 ( .A(n366), .B(n381), .C(n806), .Y(n409) );
  NAND2BXL U1518 ( .AN(n1950), .B(n362), .Y(n363) );
  NOR2XL U1519 ( .A(n1951), .B(n170), .Y(n362) );
  AOI211XL U1520 ( .A0(n1941), .A1(n1940), .B0(n1939), .C0(n1938), .Y(n1942)
         );
  NOR2XL U1521 ( .A(n1941), .B(n1940), .Y(n1938) );
  AOI211XL U1522 ( .A0(n768), .A1(n166), .B0(n200), .C0(n1937), .Y(n1939) );
  NOR2XL U1523 ( .A(n768), .B(n166), .Y(n1934) );
  INVXL U1524 ( .A(n1947), .Y(n356) );
  INVXL U1525 ( .A(n2130), .Y(n361) );
  NAND3XL U1526 ( .A(write_cntr[4]), .B(n1941), .C(n1936), .Y(n1932) );
  NAND2XL U1527 ( .A(n2131), .B(write_cntr[5]), .Y(n1923) );
  NAND2XL U1528 ( .A(n1948), .B(n1947), .Y(n2128) );
  NAND2XL U1529 ( .A(n1930), .B(n1931), .Y(n1920) );
  NOR2XL U1530 ( .A(n1913), .B(n1912), .Y(n1916) );
  INVXL U1531 ( .A(n1928), .Y(n1919) );
  INVXL U1532 ( .A(n1905), .Y(n1906) );
  NAND3XL U1533 ( .A(write_cntr[5]), .B(n1926), .C(n1941), .Y(n1918) );
  INVXL U1534 ( .A(n1902), .Y(n1904) );
  NOR2XL U1535 ( .A(n1898), .B(n1897), .Y(n1899) );
  NAND3XL U1536 ( .A(write_cntr[6]), .B(n1911), .C(n1926), .Y(n1907) );
  INVXL U1537 ( .A(n1888), .Y(n1890) );
  NAND3XL U1538 ( .A(write_cntr[7]), .B(n1895), .C(n1911), .Y(n1896) );
  NOR2XL U1539 ( .A(n1887), .B(n1886), .Y(n1881) );
  NOR2BXL U1540 ( .AN(n2144), .B(n1877), .Y(n1878) );
  NAND3XL U1541 ( .A(write_cntr[8]), .B(write_cntr[10]), .C(n1895), .Y(n1880)
         );
  NAND3XL U1542 ( .A(n202), .B(n1876), .C(n2144), .Y(n1879) );
  NAND3XL U1543 ( .A(write_cntr[9]), .B(write_cntr[11]), .C(write_cntr[10]), 
        .Y(n1876) );
  NOR2BXL U1544 ( .AN(n505), .B(n504), .Y(N91) );
  AOI21XL U1545 ( .A0(cr_read_cntr[3]), .A1(n503), .B0(n481), .Y(n504) );
  NOR2XL U1546 ( .A(cr_read_cntr[3]), .B(n479), .Y(n480) );
  NOR2BXL U1547 ( .AN(n1065), .B(n238), .Y(n1067) );
  NAND2XL U1548 ( .A(cr_read_cntr[6]), .B(n1062), .Y(n1063) );
  NAND2XL U1549 ( .A(cr_read_cntr[8]), .B(n237), .Y(n1062) );
  OAI211XL U1550 ( .A0(n2955), .A1(n1956), .B0(n2114), .C0(si_sel), .Y(n1957)
         );
  AND2XL U1551 ( .A(n1955), .B(n146), .Y(n1956) );
  NAND2XL U1552 ( .A(n2628), .B(n162), .Y(n1955) );
  INVXL U1553 ( .A(n2097), .Y(n2108) );
  AOI211XL U1554 ( .A0(n2628), .A1(n162), .B0(n68), .C0(n2955), .Y(n2097) );
  AOI21XL U1555 ( .A0(n2959), .A1(n2958), .B0(n2957), .Y(n2968) );
  AOI211XL U1556 ( .A0(N2283), .A1(n2956), .B0(n2955), .C0(n2954), .Y(n2957)
         );
  INVXL U1557 ( .A(n2960), .Y(n2961) );
  MXI2XL U1558 ( .A(n234), .B(n640), .S0(n42), .Y(n486) );
  MXI2XL U1559 ( .A(n154), .B(n632), .S0(n42), .Y(n484) );
  NAND2XL U1560 ( .A(n40), .B(\next_write_addr_w[0] ), .Y(n355) );
  NAND2XL U1561 ( .A(n40), .B(N744), .Y(n331) );
  MXI2XL U1562 ( .A(n71), .B(n137), .S0(n40), .Y(n528) );
  NAND2XL U1563 ( .A(n88), .B(n40), .Y(n346) );
  NAND2XL U1564 ( .A(n40), .B(write_addr[16]), .Y(n351) );
  NAND2XL U1565 ( .A(n42), .B(n692), .Y(n334) );
  INVXL U1566 ( .A(n624), .Y(n353) );
  NAND2XL U1567 ( .A(n2145), .B(n2945), .Y(n329) );
  NAND2XL U1568 ( .A(n40), .B(N746), .Y(n335) );
  NAND2XL U1569 ( .A(n40), .B(N747), .Y(n336) );
  NAND2XL U1570 ( .A(n40), .B(N748), .Y(n337) );
  NAND2XL U1571 ( .A(n40), .B(write_addr[9]), .Y(n328) );
  NAND2XL U1572 ( .A(write_addr[10]), .B(n40), .Y(n325) );
  MXI2XL U1573 ( .A(n659), .B(n153), .S0(n40), .Y(n490) );
  NAND2XL U1574 ( .A(n102), .B(n40), .Y(n340) );
  NAND2XL U1575 ( .A(n40), .B(n89), .Y(n343) );
  AND2XL U1576 ( .A(n620), .B(n2127), .Y(n322) );
  NAND3XL U1577 ( .A(n778), .B(n766), .C(n2113), .Y(n2127) );
  INVXL U1578 ( .A(n2121), .Y(n2123) );
  OAI211XL U1579 ( .A0(n2120), .A1(n2119), .B0(si_sel), .C0(n2118), .Y(n2124)
         );
  NAND2XL U1580 ( .A(n2644), .B(n199), .Y(n2119) );
  NOR4XL U1581 ( .A(n2117), .B(n2116), .C(n2115), .D(n2114), .Y(n2125) );
  NAND2XL U1582 ( .A(n146), .B(n2955), .Y(n2114) );
  NOR4XL U1583 ( .A(n2628), .B(n2102), .C(n73), .D(n2090), .Y(n2092) );
  NOR4BXL U1584 ( .AN(n2104), .B(n2102), .C(n199), .D(n2101), .Y(n2095) );
  INVXL U1585 ( .A(n2089), .Y(n2101) );
  NOR2XL U1586 ( .A(n2084), .B(n2085), .Y(n2083) );
  OAI2BB2XL U1587 ( .B0(work_cntr[4]), .B1(n2076), .A0N(work_cntr[4]), .A1N(
        n2076), .Y(n2091) );
  NOR2XL U1588 ( .A(n2074), .B(n2068), .Y(n2069) );
  AOI211XL U1589 ( .A0(work_cntr[5]), .A1(n2067), .B0(n2074), .C0(n2500), .Y(
        n2071) );
  INVXL U1590 ( .A(n2085), .Y(n2077) );
  INVXL U1591 ( .A(n2073), .Y(n2067) );
  AOI211XL U1592 ( .A0(n2148), .A1(n2066), .B0(n2075), .C0(n2060), .Y(n2065)
         );
  NAND2XL U1593 ( .A(n2062), .B(n2061), .Y(n2054) );
  INVXL U1594 ( .A(n2063), .Y(n2057) );
  NAND3XL U1595 ( .A(n2058), .B(n2072), .C(n2061), .Y(n2063) );
  INVXL U1596 ( .A(n2060), .Y(n2072) );
  NAND2BXL U1597 ( .AN(n2039), .B(n2038), .Y(n2044) );
  INVXL U1598 ( .A(n2037), .Y(n2045) );
  AOI211XL U1599 ( .A0(n110), .A1(n2037), .B0(n2028), .C0(n2033), .Y(n2029) );
  NOR2BXL U1600 ( .AN(n2039), .B(n2031), .Y(n2022) );
  AOI32XL U1601 ( .A0(n2038), .A1(n2021), .A2(n2026), .B0(n2039), .B1(n2021), 
        .Y(n2024) );
  XNOR2XL U1602 ( .A(n113), .B(n2020), .Y(n2025) );
  INVXL U1603 ( .A(n2021), .Y(n2031) );
  AND2XL U1604 ( .A(n2026), .B(n2038), .Y(n2032) );
  INVXL U1605 ( .A(n2028), .Y(n2038) );
  NOR2XL U1606 ( .A(n2018), .B(n2017), .Y(n2015) );
  NAND3XL U1607 ( .A(n2012), .B(n2010), .C(n2018), .Y(n2011) );
  NAND3XL U1608 ( .A(n113), .B(n2019), .C(n2016), .Y(n2010) );
  NAND2XL U1609 ( .A(n2009), .B(n2008), .Y(n2019) );
  INVXL U1610 ( .A(n2017), .Y(n2012) );
  NOR2BXL U1611 ( .AN(n2005), .B(n2004), .Y(n2023) );
  AOI211XL U1612 ( .A0(n2009), .A1(n2005), .B0(n1999), .C0(n2004), .Y(n2001)
         );
  INVXL U1613 ( .A(n2006), .Y(n1999) );
  NOR2XL U1614 ( .A(work_cntr[11]), .B(n2541), .Y(n1996) );
  INVXL U1615 ( .A(n1989), .Y(n2003) );
  INVXL U1616 ( .A(n2007), .Y(n1990) );
  NAND2XL U1617 ( .A(n1984), .B(n1983), .Y(n1985) );
  NAND2XL U1618 ( .A(n1982), .B(n1981), .Y(n1986) );
  NAND2BXL U1619 ( .AN(n1980), .B(n1979), .Y(n1981) );
  NOR2XL U1620 ( .A(n1978), .B(n1977), .Y(n1975) );
  NOR3XL U1621 ( .A(n1978), .B(n1980), .C(n1979), .Y(n1976) );
  NAND2XL U1622 ( .A(n1979), .B(n1980), .Y(n1977) );
  NAND2XL U1623 ( .A(n1982), .B(n1974), .Y(n1980) );
  INVXL U1624 ( .A(n1973), .Y(n1978) );
  XOR2XL U1625 ( .A(n1969), .B(n1968), .Y(n1970) );
  NAND4XL U1626 ( .A(n1979), .B(n1973), .C(n1982), .D(n1968), .Y(n1964) );
  INVXL U1627 ( .A(n1974), .Y(n1968) );
  NAND2XL U1628 ( .A(n2014), .B(n1960), .Y(n1961) );
  INVXL U1629 ( .A(n2148), .Y(n2068) );
  AOI222XL U1630 ( .A0(n254), .A1(\C168/DATA3_0 ), .B0(n779), .B1(
        global_cntr[0]), .C0(n759), .C1(N1667), .Y(\im_a[0]_BAR ) );
  MXI2XL U1631 ( .A(n151), .B(n2971), .S0(read_cntr[0]), .Y(n521) );
  AOI211XL U1632 ( .A0(n245), .A1(n358), .B0(n359), .C0(n41), .Y(n501) );
  NAND2XL U1633 ( .A(n69), .B(N1453), .Y(n358) );
  AOI211XL U1634 ( .A0(n240), .A1(n2934), .B0(n2935), .C0(n41), .Y(n499) );
  AOI211XL U1635 ( .A0(n2936), .A1(n241), .B0(n2937), .C0(n41), .Y(n498) );
  INVXL U1636 ( .A(n2938), .Y(n497) );
  OAI211XL U1637 ( .A0(n2937), .A1(cr_read_cntr[5]), .B0(n2939), .C0(n257), 
        .Y(n2938) );
  AOI211XL U1638 ( .A0(n2939), .A1(n242), .B0(n2940), .C0(n41), .Y(n496) );
  AOI211XL U1639 ( .A0(n2941), .A1(n237), .B0(n2943), .C0(n41), .Y(n495) );
  AOI211XL U1640 ( .A0(cr_read_cntr[8]), .A1(n2943), .B0(n41), .C0(n2942), .Y(
        n494) );
  NOR2XL U1641 ( .A(cr_read_cntr[8]), .B(n2943), .Y(n2942) );
  INVXL U1642 ( .A(n2940), .Y(n2941) );
  INVXL U1643 ( .A(n2935), .Y(n2936) );
  NAND2XL U1644 ( .A(n359), .B(N1455), .Y(n2934) );
  NOR2XL U1645 ( .A(n2916), .B(n2917), .Y(n2915) );
  INVXL U1646 ( .A(n2914), .Y(n2917) );
  AOI211XL U1647 ( .A0(n2912), .A1(n2911), .B0(n2910), .C0(n2909), .Y(n2920)
         );
  NOR2XL U1648 ( .A(n2912), .B(n2911), .Y(n2909) );
  NAND3XL U1649 ( .A(n2908), .B(n2907), .C(n2906), .Y(n2910) );
  AOI211XL U1650 ( .A0(n2905), .A1(n2904), .B0(n2903), .C0(n2902), .Y(n2906)
         );
  NOR3XL U1651 ( .A(n2905), .B(n2901), .C(n2904), .Y(n2902) );
  NOR3XL U1652 ( .A(n2900), .B(n772), .C(n2899), .Y(n2907) );
  NAND2XL U1653 ( .A(n2897), .B(n2913), .Y(n2914) );
  INVXL U1654 ( .A(n2892), .Y(n2895) );
  NAND2BXL U1655 ( .AN(n2905), .B(n2904), .Y(n2896) );
  NAND2XL U1656 ( .A(n2878), .B(n2888), .Y(n2881) );
  NAND3XL U1657 ( .A(n2882), .B(n2884), .C(n2877), .Y(n2888) );
  NAND3XL U1658 ( .A(n2874), .B(n2871), .C(n2870), .Y(n2872) );
  NOR4BXL U1659 ( .AN(n2869), .B(next_work_cntr[2]), .C(n2868), .D(n2867), .Y(
        n2871) );
  NAND2XL U1660 ( .A(n2870), .B(n2876), .Y(n2878) );
  NAND2XL U1661 ( .A(n2857), .B(n2856), .Y(n2854) );
  INVXL U1662 ( .A(n2849), .Y(n2850) );
  NAND2BXL U1663 ( .AN(n2848), .B(n2876), .Y(n2856) );
  INVXL U1664 ( .A(n2843), .Y(n2846) );
  NOR2XL U1665 ( .A(n2838), .B(n2837), .Y(n2840) );
  NAND3XL U1666 ( .A(n2870), .B(n2834), .C(n2869), .Y(n2842) );
  NAND2XL U1667 ( .A(n2831), .B(n2882), .Y(n2848) );
  INVXL U1668 ( .A(n2834), .Y(n2868) );
  INVXL U1669 ( .A(n2880), .Y(n2889) );
  NAND3XL U1670 ( .A(n2823), .B(n2825), .C(n2832), .Y(n2824) );
  NAND2XL U1671 ( .A(n2833), .B(n2862), .Y(n2823) );
  NAND2XL U1672 ( .A(n2831), .B(n2851), .Y(n2827) );
  INVXL U1673 ( .A(n2821), .Y(n2833) );
  NAND2XL U1674 ( .A(n2844), .B(n2843), .Y(n2819) );
  INVXL U1675 ( .A(n2815), .Y(n2818) );
  NAND2XL U1676 ( .A(n2839), .B(n2845), .Y(n2844) );
  NAND4XL U1677 ( .A(n2808), .B(n2807), .C(n2831), .D(n2820), .Y(n2809) );
  INVXL U1678 ( .A(n2802), .Y(n2804) );
  NAND3XL U1679 ( .A(n2801), .B(n2798), .C(n2800), .Y(n2799) );
  NAND2XL U1680 ( .A(n2802), .B(n2803), .Y(n2798) );
  INVXL U1681 ( .A(n2858), .Y(n2806) );
  INVXL U1682 ( .A(n2791), .Y(n2793) );
  NAND2XL U1683 ( .A(n2817), .B(n2790), .Y(n2816) );
  NAND4XL U1684 ( .A(n2808), .B(n2858), .C(n2789), .D(n2802), .Y(n2790) );
  INVXL U1685 ( .A(n2782), .Y(n2784) );
  NOR2XL U1686 ( .A(n2813), .B(n2812), .Y(n2780) );
  INVXL U1687 ( .A(n2767), .Y(n2770) );
  NAND2XL U1688 ( .A(n2794), .B(n2779), .Y(n2792) );
  NAND3XL U1689 ( .A(n2778), .B(n2788), .C(n2766), .Y(n2779) );
  NOR4XL U1690 ( .A(next_work_cntr[5]), .B(n78), .C(n2822), .D(n2772), .Y(
        n2766) );
  AND2XL U1691 ( .A(n2811), .B(n2786), .Y(n2778) );
  NAND2XL U1692 ( .A(n2752), .B(n2807), .Y(n2772) );
  INVXL U1693 ( .A(n2774), .Y(n2754) );
  NAND2XL U1694 ( .A(n2768), .B(n2767), .Y(n2750) );
  INVXL U1695 ( .A(n2742), .Y(n2745) );
  NAND2XL U1696 ( .A(n2728), .B(n2736), .Y(n2757) );
  INVXL U1697 ( .A(n2776), .Y(n2752) );
  NAND2XL U1698 ( .A(n2786), .B(n80), .Y(n2756) );
  OAI2BB2XL U1699 ( .B0(n2725), .B1(n2724), .A0N(n2725), .A1N(n2724), .Y(n2783) );
  NAND2XL U1700 ( .A(n2743), .B(n2742), .Y(n2734) );
  NAND2XL U1701 ( .A(n2744), .B(n2739), .Y(n2743) );
  NAND2XL U1702 ( .A(n2761), .B(n2758), .Y(n2741) );
  INVXL U1703 ( .A(n2725), .Y(n2720) );
  INVXL U1704 ( .A(n2704), .Y(n2706) );
  INVXL U1705 ( .A(n2749), .Y(n2735) );
  NAND2BXL U1706 ( .AN(n2702), .B(n2698), .Y(n2699) );
  AND2XL U1707 ( .A(n2712), .B(n2709), .Y(n2729) );
  AND2XL U1708 ( .A(n2727), .B(n2722), .Y(n2709) );
  NAND2XL U1709 ( .A(n2731), .B(n2732), .Y(n2704) );
  INVXL U1710 ( .A(n2696), .Y(n2701) );
  INVXL U1711 ( .A(n2692), .Y(n2694) );
  NAND2XL U1712 ( .A(n2718), .B(n2696), .Y(n2717) );
  NAND4BXL U1713 ( .AN(n2691), .B(n2690), .C(n2712), .D(n2689), .Y(n2696) );
  NOR3XL U1714 ( .A(n2703), .B(n2716), .C(n2700), .Y(n2689) );
  NAND3XL U1715 ( .A(n2728), .B(n2727), .C(n2731), .Y(n2716) );
  INVXL U1716 ( .A(n2710), .Y(n2676) );
  INVXL U1717 ( .A(n2698), .Y(n2703) );
  INVXL U1718 ( .A(n2672), .Y(n2674) );
  INVXL U1719 ( .A(n2669), .Y(n2682) );
  NOR3XL U1720 ( .A(next_work_cntr[15]), .B(next_work_cntr[16]), .C(n2662), 
        .Y(n2665) );
  NAND2XL U1721 ( .A(n2688), .B(n2687), .Y(n2668) );
  INVXL U1722 ( .A(n2675), .Y(n2662) );
  NAND2XL U1723 ( .A(n2714), .B(n2715), .Y(n2672) );
  NAND2XL U1724 ( .A(next_work_cntr[18]), .B(n2663), .Y(n2692) );
  NAND3XL U1725 ( .A(next_work_cntr[18]), .B(n2657), .C(next_work_cntr[19]), 
        .Y(n2663) );
  NAND2XL U1726 ( .A(n2714), .B(n2658), .Y(n2691) );
  INVXL U1727 ( .A(n2707), .Y(n2658) );
  NAND2XL U1728 ( .A(n2678), .B(n2650), .Y(n2669) );
  NAND2XL U1729 ( .A(n2657), .B(n2648), .Y(n2655) );
  OR3XL U1730 ( .A(n2680), .B(next_work_cntr[14]), .C(next_work_cntr[10]), .Y(
        n2651) );
  OAI211XL U1731 ( .A0(n2647), .A1(n2646), .B0(n2962), .C0(n2645), .Y(n2922)
         );
  XNOR2XL U1732 ( .A(n2641), .B(n2640), .Y(n2642) );
  AOI21XL U1733 ( .A0(n2643), .A1(N2282), .B0(N205), .Y(n2641) );
  NAND3XL U1734 ( .A(n2630), .B(n2632), .C(n2635), .Y(n2631) );
  AND2XL U1735 ( .A(n2632), .B(n2635), .Y(n2622) );
  INVXL U1736 ( .A(n2620), .Y(n2627) );
  INVXL U1737 ( .A(n2626), .Y(n2616) );
  INVXL U1738 ( .A(n2614), .Y(n2612) );
  NAND3XL U1739 ( .A(n2607), .B(n2604), .C(n2606), .Y(n2605) );
  AND2XL U1740 ( .A(n2613), .B(n2615), .Y(n2619) );
  NOR2XL U1741 ( .A(work_cntr[4]), .B(n2608), .Y(n2592) );
  INVXL U1742 ( .A(n2602), .Y(n2603) );
  NAND3XL U1743 ( .A(n2596), .B(n2597), .C(n2593), .Y(n2604) );
  NAND3XL U1744 ( .A(n2595), .B(n2594), .C(n2590), .Y(n2593) );
  INVXL U1745 ( .A(n2589), .Y(n2595) );
  INVXL U1746 ( .A(n2585), .Y(n2583) );
  INVXL U1747 ( .A(n2581), .Y(n2574) );
  INVXL U1748 ( .A(n2571), .Y(n2572) );
  NOR3XL U1749 ( .A(n2556), .B(n2562), .C(n2564), .Y(n2557) );
  INVXL U1750 ( .A(n2565), .Y(n2556) );
  NOR3XL U1751 ( .A(n2538), .B(n2542), .C(n2544), .Y(n2539) );
  NAND2XL U1752 ( .A(n2529), .B(n2528), .Y(n2533) );
  INVXL U1753 ( .A(n2524), .Y(n2527) );
  NOR2XL U1754 ( .A(n2542), .B(n2535), .Y(n2536) );
  INVXL U1755 ( .A(n2525), .Y(n2517) );
  NAND2XL U1756 ( .A(n2513), .B(n2512), .Y(n2524) );
  NAND2XL U1757 ( .A(n2514), .B(n2526), .Y(n2519) );
  INVXL U1758 ( .A(n2510), .Y(n2511) );
  NAND2BXL U1759 ( .AN(n2512), .B(n2510), .Y(n2514) );
  NOR2XL U1760 ( .A(n2508), .B(work_cntr[19]), .Y(n2507) );
  INVXL U1761 ( .A(n2520), .Y(n2531) );
  NAND2XL U1762 ( .A(n2503), .B(n2502), .Y(n2504) );
  INVXL U1763 ( .A(n2521), .Y(n2503) );
  NAND2XL U1764 ( .A(n2492), .B(n2490), .Y(n2491) );
  NOR2BXL U1765 ( .AN(n2488), .B(n2487), .Y(n2489) );
  NOR2XL U1766 ( .A(n2493), .B(n2492), .Y(n2483) );
  NAND2XL U1767 ( .A(n2494), .B(n2484), .Y(n2488) );
  INVXL U1768 ( .A(n2477), .Y(n2474) );
  INVXL U1769 ( .A(n2473), .Y(n2479) );
  INVXL U1770 ( .A(n2485), .Y(n2494) );
  NOR2XL U1771 ( .A(n2476), .B(n2473), .Y(n2471) );
  NAND2XL U1772 ( .A(n2472), .B(n2477), .Y(n2481) );
  NAND2XL U1773 ( .A(n2467), .B(n2469), .Y(n2477) );
  NAND2BXL U1774 ( .AN(n59), .B(n2465), .Y(n2469) );
  NAND2XL U1775 ( .A(n2461), .B(n2460), .Y(n2465) );
  NAND2XL U1776 ( .A(n59), .B(n2459), .Y(n2467) );
  NAND2XL U1777 ( .A(n44), .B(n2470), .Y(n2459) );
  NAND2XL U1778 ( .A(n2456), .B(n2454), .Y(n2455) );
  NOR2XL U1779 ( .A(n2457), .B(n2456), .Y(n2451) );
  NAND2XL U1780 ( .A(n2452), .B(n2458), .Y(n2460) );
  NAND2XL U1781 ( .A(n2447), .B(n2449), .Y(n2458) );
  NAND2BXL U1782 ( .AN(n2446), .B(n2445), .Y(n2449) );
  NAND2XL U1783 ( .A(n2441), .B(n2440), .Y(n2445) );
  NAND2XL U1784 ( .A(n2446), .B(n2439), .Y(n2447) );
  NAND2XL U1785 ( .A(n45), .B(n2450), .Y(n2439) );
  NAND2XL U1786 ( .A(n2436), .B(n2434), .Y(n2435) );
  NOR2XL U1787 ( .A(n2437), .B(n2436), .Y(n2432) );
  NAND2XL U1788 ( .A(n53), .B(n2438), .Y(n2440) );
  NAND2BXL U1789 ( .AN(n2426), .B(n2425), .Y(n2429) );
  NAND2XL U1790 ( .A(n2421), .B(n2420), .Y(n2425) );
  NAND2XL U1791 ( .A(n2426), .B(n2419), .Y(n2427) );
  NAND2XL U1792 ( .A(n2424), .B(n2430), .Y(n2419) );
  NAND2XL U1793 ( .A(n2416), .B(n2414), .Y(n2415) );
  NOR2XL U1794 ( .A(n2417), .B(n2416), .Y(n2412) );
  INVXL U1795 ( .A(n2413), .Y(n2417) );
  NAND2XL U1796 ( .A(n2411), .B(n2418), .Y(n2420) );
  NAND2BXL U1797 ( .AN(n2406), .B(n2405), .Y(n2409) );
  NAND2XL U1798 ( .A(n2401), .B(n2400), .Y(n2405) );
  NAND2XL U1799 ( .A(n2406), .B(n2399), .Y(n2407) );
  NAND2XL U1800 ( .A(n2404), .B(n2410), .Y(n2399) );
  NAND2XL U1801 ( .A(n2397), .B(n2395), .Y(n2396) );
  NOR2XL U1802 ( .A(n2649), .B(n2397), .Y(n2392) );
  NAND2XL U1803 ( .A(n49), .B(n2398), .Y(n2400) );
  NAND2BXL U1804 ( .AN(n2388), .B(n2387), .Y(n2391) );
  NAND2XL U1805 ( .A(n2383), .B(n2382), .Y(n2387) );
  NAND2XL U1806 ( .A(n2388), .B(n2381), .Y(n2389) );
  NAND2XL U1807 ( .A(n2386), .B(n2671), .Y(n2381) );
  NAND2XL U1808 ( .A(n2378), .B(n2376), .Y(n2377) );
  NOR2XL U1809 ( .A(n2379), .B(n2378), .Y(n2373) );
  NAND2XL U1810 ( .A(n50), .B(n2380), .Y(n2382) );
  NAND2BXL U1811 ( .AN(n2368), .B(n2367), .Y(n2371) );
  NAND2XL U1812 ( .A(n2364), .B(n2363), .Y(n2367) );
  NAND2XL U1813 ( .A(n2362), .B(n2368), .Y(n2369) );
  NAND2XL U1814 ( .A(n2359), .B(n2357), .Y(n2358) );
  NAND2XL U1815 ( .A(n2366), .B(n2372), .Y(n2362) );
  NOR2XL U1816 ( .A(n2360), .B(n2359), .Y(n2354) );
  NAND2XL U1817 ( .A(n2355), .B(n2361), .Y(n2363) );
  NAND2XL U1818 ( .A(n2349), .B(n2348), .Y(n2352) );
  NAND2XL U1819 ( .A(n2345), .B(n2344), .Y(n2348) );
  NOR2XL U1820 ( .A(n2660), .B(n2342), .Y(n2343) );
  INVXL U1821 ( .A(n2342), .Y(n2347) );
  NAND2XL U1822 ( .A(n2335), .B(n2334), .Y(n2345) );
  NAND2XL U1823 ( .A(n2341), .B(n2336), .Y(n2334) );
  NAND2BXL U1824 ( .AN(n2335), .B(n2338), .Y(n2344) );
  NAND2XL U1825 ( .A(n2331), .B(n2330), .Y(n2338) );
  NOR2BXL U1826 ( .AN(n2329), .B(n2333), .Y(n2331) );
  NAND2XL U1827 ( .A(work_cntr[19]), .B(n2326), .Y(n2327) );
  NOR2XL U1828 ( .A(n2333), .B(n2332), .Y(n2328) );
  INVXL U1829 ( .A(n2321), .Y(n2323) );
  AOI31XL U1830 ( .A0(n2320), .A1(n2319), .A2(n2318), .B0(n2317), .Y(n2325) );
  NOR4XL U1831 ( .A(n2316), .B(n2315), .C(n2314), .D(n2313), .Y(n2317) );
  NAND4XL U1832 ( .A(n2671), .B(n2356), .C(n2336), .D(n2375), .Y(n2314) );
  NAND4XL U1833 ( .A(n2311), .B(n2430), .C(n2372), .D(n2353), .Y(n2315) );
  NOR4XL U1834 ( .A(n2402), .B(n2457), .C(n2310), .D(n2309), .Y(n2311) );
  NAND4XL U1835 ( .A(n2450), .B(n2394), .C(n2413), .D(n2433), .Y(n2316) );
  INVXL U1836 ( .A(n2437), .Y(n2433) );
  NAND2XL U1837 ( .A(n2308), .B(n2654), .Y(n2318) );
  NAND3XL U1838 ( .A(n2307), .B(n2306), .C(n2305), .Y(n2304) );
  NAND3XL U1839 ( .A(n2300), .B(n2297), .C(n2299), .Y(n2298) );
  NAND2XL U1840 ( .A(n2296), .B(n2301), .Y(n2297) );
  OAI211XL U1841 ( .A0(n2300), .A1(n2295), .B0(n2293), .C0(n2296), .Y(n2292)
         );
  INVXL U1842 ( .A(n2303), .Y(n2295) );
  NAND2XL U1843 ( .A(n199), .B(n257), .Y(n2303) );
  INVXL U1844 ( .A(n2294), .Y(n2296) );
  INVXL U1845 ( .A(n2291), .Y(n2287) );
  OAI211XL U1846 ( .A0(n2291), .A1(n2284), .B0(n2279), .C0(n2286), .Y(n2283)
         );
  OAI211XL U1847 ( .A0(n2276), .A1(n2271), .B0(n2272), .C0(n2266), .Y(n2268)
         );
  NAND2XL U1848 ( .A(n2265), .B(n2264), .Y(n2272) );
  NAND2BXL U1849 ( .AN(n2263), .B(n2262), .Y(n2264) );
  INVXL U1850 ( .A(n2275), .Y(n2269) );
  INVXL U1851 ( .A(n2261), .Y(n2266) );
  NAND2XL U1852 ( .A(n2249), .B(n2258), .Y(n2248) );
  NAND2XL U1853 ( .A(n2245), .B(n2244), .Y(n2258) );
  NAND2XL U1854 ( .A(n2241), .B(n2240), .Y(n2242) );
  NAND2XL U1855 ( .A(n2247), .B(n2246), .Y(n2240) );
  AND2XL U1856 ( .A(n2236), .B(n2235), .Y(n2243) );
  AOI211XL U1857 ( .A0(n2239), .A1(n2241), .B0(n2230), .C0(n2237), .Y(n2232)
         );
  INVXL U1858 ( .A(n2235), .Y(n2230) );
  OAI211XL U1859 ( .A0(n2222), .A1(n2221), .B0(n2224), .C0(n2225), .Y(n2223)
         );
  INVXL U1860 ( .A(n2231), .Y(n2221) );
  NAND3XL U1861 ( .A(n2236), .B(n2235), .C(n2228), .Y(n2219) );
  NAND2XL U1862 ( .A(n2216), .B(n2215), .Y(n2235) );
  NAND2BXL U1863 ( .AN(n2214), .B(n2220), .Y(n2233) );
  INVXL U1864 ( .A(n2211), .Y(n2215) );
  INVXL U1865 ( .A(n2200), .Y(n2201) );
  NAND2XL U1866 ( .A(n2204), .B(n2199), .Y(n2205) );
  INVXL U1867 ( .A(n2213), .Y(n2197) );
  NOR2XL U1868 ( .A(next_work_cntr[11]), .B(n2217), .Y(n2194) );
  INVXL U1869 ( .A(n2202), .Y(n2210) );
  INVXL U1870 ( .A(n2181), .Y(n2183) );
  INVXL U1871 ( .A(n2189), .Y(n2206) );
  INVXL U1872 ( .A(n2191), .Y(n2186) );
  AOI211XL U1873 ( .A0(n2176), .A1(n2175), .B0(n2182), .C0(n2174), .Y(n2177)
         );
  NOR2XL U1874 ( .A(n2173), .B(n2176), .Y(n2174) );
  INVXL U1875 ( .A(n2171), .Y(n2175) );
  NAND2XL U1876 ( .A(n2173), .B(n2168), .Y(n2171) );
  OAI211XL U1877 ( .A0(n2163), .A1(n2162), .B0(n2173), .C0(n2166), .Y(n2164)
         );
  AND3XL U1878 ( .A(n2163), .B(n2162), .C(n2173), .Y(n2165) );
  NAND2XL U1879 ( .A(n2160), .B(n2163), .Y(n2168) );
  NOR2XL U1880 ( .A(next_work_cntr[15]), .B(n2167), .Y(n2159) );
  NOR2BXL U1881 ( .AN(n2163), .B(n2160), .Y(n2161) );
  NAND2BXL U1882 ( .AN(n2167), .B(n2156), .Y(n2158) );
  INVXL U1883 ( .A(n2664), .Y(next_work_cntr[17]) );
  INVXL U1884 ( .A(n2155), .Y(n2308) );
  NAND2XL U1885 ( .A(n2157), .B(n2648), .Y(n2155) );
  INVXL U1886 ( .A(n2336), .Y(n2337) );
  INVXL U1887 ( .A(n1033), .Y(n1032) );
  NAND2XL U1888 ( .A(work_cntr[16]), .B(n1034), .Y(n1033) );
  INVXL U1889 ( .A(n2450), .Y(n2442) );
  INVXL U1890 ( .A(n2733), .Y(next_work_cntr[7]) );
  INVXL U1891 ( .A(n2430), .Y(n2422) );
  NAND2XL U1892 ( .A(n129), .B(n1044), .Y(n1043) );
  AOI222XL U1893 ( .A0(n254), .A1(\C168/DATA3_19 ), .B0(global_cntr[19]), .B1(
        n779), .C0(n759), .C1(N1686), .Y(\im_a[19]_BAR ) );
  INVXL U1894 ( .A(n2110), .Y(n2112) );
  NOR2XL U1895 ( .A(n2113), .B(sftr_n[1]), .Y(n721) );
  NOR2BXL U1896 ( .AN(curr_photo_addr[19]), .B(n718), .Y(\C1/Z_19 ) );
  AOI211XL U1897 ( .A0(write_addr[17]), .A1(n649), .B0(n626), .C0(n625), .Y(
        n627) );
  NOR2XL U1898 ( .A(n632), .B(n703), .Y(n626) );
  AOI211XL U1899 ( .A0(n2145), .A1(n707), .B0(n706), .C0(n705), .Y(n708) );
  NOR2XL U1900 ( .A(n711), .B(n703), .Y(n706) );
  OAI211XL U1901 ( .A0(n612), .A1(n71), .B0(n611), .C0(n610), .Y(\C169/Z_1 )
         );
  NAND2XL U1902 ( .A(N743), .B(n609), .Y(n610) );
  AOI22XL U1903 ( .A0(N622), .A1(n252), .B0(N743), .B1(n253), .Y(n611) );
  AOI211XL U1904 ( .A0(n1087), .A1(n1086), .B0(n1431), .C0(n1085), .Y(n1159)
         );
  NOR2XL U1905 ( .A(\next_write_addr_w[0] ), .B(n1087), .Y(n1085) );
  OAI211XL U1906 ( .A0(n1283), .A1(n1155), .B0(n251), .C0(n1291), .Y(n1156) );
  NAND2XL U1907 ( .A(n1369), .B(n1084), .Y(n1157) );
  INVXL U1908 ( .A(n1084), .Y(n354) );
  NAND2XL U1909 ( .A(n781), .B(n1072), .Y(n1084) );
  OAI211XL U1910 ( .A0(n618), .A1(n173), .B0(n617), .C0(n616), .Y(\C169/Z_0 )
         );
  NAND2XL U1911 ( .A(n2145), .B(n615), .Y(n616) );
  AOI22XL U1912 ( .A0(n173), .A1(n252), .B0(N742), .B1(n253), .Y(n617) );
  NOR2BXL U1913 ( .AN(curr_photo_addr[0]), .B(n718), .Y(n761) );
  AOI211XL U1914 ( .A0(n701), .A1(n2145), .B0(n700), .C0(n699), .Y(n702) );
  NOR2XL U1915 ( .A(n71), .B(n712), .Y(n700) );
  OAI211XL U1916 ( .A0(n618), .A1(n211), .B0(n608), .C0(n607), .Y(\C169/Z_2 )
         );
  NAND2XL U1917 ( .A(n615), .B(n696), .Y(n607) );
  AOI22XL U1918 ( .A0(N623), .A1(n252), .B0(N744), .B1(n253), .Y(n608) );
  AOI211XL U1919 ( .A0(n707), .A1(n696), .B0(n695), .C0(n694), .Y(n697) );
  NOR2XL U1920 ( .A(n71), .B(n703), .Y(n695) );
  AOI211XL U1921 ( .A0(n776), .A1(N743), .B0(n1417), .C0(n330), .Y(n698) );
  AOI211XL U1922 ( .A0(n173), .A1(n137), .B0(n1431), .C0(n1416), .Y(n330) );
  AOI211XL U1923 ( .A0(n1415), .A1(n1414), .B0(n1428), .C0(n1413), .Y(n1417)
         );
  NOR2XL U1924 ( .A(n1415), .B(n1414), .Y(n1413) );
  OAI211XL U1925 ( .A0(n618), .A1(n167), .B0(n606), .C0(n605), .Y(\C169/Z_3 )
         );
  NAND2XL U1926 ( .A(n615), .B(n692), .Y(n605) );
  AOI22XL U1927 ( .A0(N624), .A1(n252), .B0(N745), .B1(n253), .Y(n606) );
  AOI211XL U1928 ( .A0(n707), .A1(n692), .B0(n691), .C0(n690), .Y(n693) );
  NOR2XL U1929 ( .A(n689), .B(n703), .Y(n691) );
  INVXL U1930 ( .A(n696), .Y(n689) );
  OAI211XL U1931 ( .A0(n612), .A1(n685), .B0(n604), .C0(n603), .Y(\C169/Z_4 )
         );
  NAND2XL U1932 ( .A(N746), .B(n609), .Y(n603) );
  AOI22XL U1933 ( .A0(N625), .A1(n252), .B0(N746), .B1(n253), .Y(n604) );
  NOR2BXL U1934 ( .AN(curr_photo_addr[5]), .B(n718), .Y(\C1/Z_5 ) );
  AOI211XL U1935 ( .A0(n701), .A1(n692), .B0(n687), .C0(n686), .Y(n688) );
  NOR2XL U1936 ( .A(n685), .B(n712), .Y(n687) );
  AOI21XL U1937 ( .A0(n776), .A1(N745), .B0(n332), .Y(n333) );
  AOI211XL U1938 ( .A0(n1424), .A1(n167), .B0(n1431), .C0(n1423), .Y(n332) );
  OAI211XL U1939 ( .A0(n618), .A1(n136), .B0(n602), .C0(n601), .Y(\C169/Z_5 )
         );
  NAND2XL U1940 ( .A(n615), .B(n683), .Y(n601) );
  AOI22XL U1941 ( .A0(N626), .A1(n252), .B0(N747), .B1(n253), .Y(n602) );
  NOR2BXL U1942 ( .AN(curr_photo_addr[6]), .B(n718), .Y(\C1/Z_6 ) );
  AOI211XL U1943 ( .A0(n707), .A1(n683), .B0(n682), .C0(n681), .Y(n684) );
  NOR2XL U1944 ( .A(n685), .B(n703), .Y(n682) );
  OAI211XL U1945 ( .A0(n612), .A1(n677), .B0(n600), .C0(n599), .Y(\C169/Z_6 )
         );
  NAND2XL U1946 ( .A(N748), .B(n609), .Y(n599) );
  AOI22XL U1947 ( .A0(N627), .A1(n252), .B0(N748), .B1(n253), .Y(n600) );
  AOI211XL U1948 ( .A0(n701), .A1(n683), .B0(n679), .C0(n678), .Y(n680) );
  NOR2XL U1949 ( .A(n677), .B(n712), .Y(n679) );
  OAI211XL U1950 ( .A0(n612), .A1(n668), .B0(n596), .C0(n595), .Y(\C169/Z_7 )
         );
  NOR2XL U1951 ( .A(n171), .B(n597), .Y(n594) );
  AOI22XL U1952 ( .A0(N628), .A1(n252), .B0(n233), .B1(n253), .Y(n596) );
  NOR2BXL U1953 ( .AN(curr_photo_addr[8]), .B(n718), .Y(\C1/Z_8 ) );
  AOI211XL U1954 ( .A0(n707), .A1(n675), .B0(n674), .C0(n673), .Y(n676) );
  NOR2XL U1955 ( .A(n677), .B(n703), .Y(n674) );
  OAI211XL U1956 ( .A0(n664), .A1(n612), .B0(n592), .C0(n591), .Y(\C169/Z_8 )
         );
  NAND2XL U1957 ( .A(write_addr[10]), .B(n593), .Y(n591) );
  NAND2XL U1958 ( .A(n598), .B(n1719), .Y(n593) );
  AOI211XL U1959 ( .A0(N629), .A1(n252), .B0(n590), .C0(n589), .Y(n592) );
  NOR4XL U1960 ( .A(n597), .B(write_addr[10]), .C(n171), .D(n233), .Y(n589) );
  AND2XL U1961 ( .A(N750), .B(n253), .Y(n590) );
  NOR2BXL U1962 ( .AN(curr_photo_addr[9]), .B(n718), .Y(\C1/Z_9 ) );
  INVXL U1963 ( .A(n668), .Y(n671) );
  AOI211XL U1964 ( .A0(N630), .A1(n252), .B0(n587), .C0(n586), .Y(n588) );
  AOI211XL U1965 ( .A0(n1720), .A1(n153), .B0(n597), .C0(n770), .Y(n585) );
  NOR2XL U1966 ( .A(n598), .B(n153), .Y(n587) );
  NOR2BXL U1967 ( .AN(curr_photo_addr[10]), .B(n718), .Y(\C1/Z_10 ) );
  AOI211XL U1968 ( .A0(n701), .A1(n675), .B0(n666), .C0(n665), .Y(n667) );
  NOR2XL U1969 ( .A(n664), .B(n712), .Y(n666) );
  AOI211XL U1970 ( .A0(n1404), .A1(n1369), .B0(n2926), .C0(n1317), .Y(n1318)
         );
  OAI211XL U1971 ( .A0(n654), .A1(n612), .B0(n584), .C0(n583), .Y(\C169/Z_10 )
         );
  NOR2XL U1972 ( .A(n597), .B(n580), .Y(n582) );
  INVXL U1973 ( .A(n770), .Y(n580) );
  AOI22XL U1974 ( .A0(N631), .A1(n252), .B0(N752), .B1(n253), .Y(n584) );
  AOI211XL U1975 ( .A0(n707), .A1(n662), .B0(n661), .C0(n660), .Y(n663) );
  NOR2XL U1976 ( .A(n668), .B(n703), .Y(n661) );
  NAND2XL U1977 ( .A(n776), .B(write_addr[9]), .Y(n326) );
  AOI211XL U1978 ( .A0(n1369), .A1(n1370), .B0(n1368), .C0(n1398), .Y(n1371)
         );
  INVXL U1979 ( .A(n659), .Y(n662) );
  OAI211XL U1980 ( .A0(n612), .A1(n648), .B0(n579), .C0(n578), .Y(\C169/Z_11 )
         );
  NAND2XL U1981 ( .A(n89), .B(n581), .Y(n578) );
  AOI211XL U1982 ( .A0(N632), .A1(n252), .B0(n577), .C0(n576), .Y(n579) );
  AND2XL U1983 ( .A(n770), .B(n102), .Y(n1714) );
  AND2XL U1984 ( .A(N753), .B(n253), .Y(n577) );
  NOR2BXL U1985 ( .AN(curr_photo_addr[12]), .B(n718), .Y(\C1/Z_12 ) );
  AOI211XL U1986 ( .A0(n707), .A1(n657), .B0(n656), .C0(n655), .Y(n658) );
  NOR2XL U1987 ( .A(n664), .B(n703), .Y(n656) );
  NAND2XL U1988 ( .A(n776), .B(write_addr[10]), .Y(n323) );
  AOI211XL U1989 ( .A0(n1314), .A1(n1315), .B0(n1362), .C0(n1398), .Y(n1316)
         );
  NOR2XL U1990 ( .A(n233), .B(n1366), .Y(n1313) );
  INVXL U1991 ( .A(n1368), .Y(n1314) );
  INVXL U1992 ( .A(n654), .Y(n657) );
  OAI211XL U1993 ( .A0(n644), .A1(n612), .B0(n575), .C0(n574), .Y(\C169/Z_12 )
         );
  INVXL U1994 ( .A(n571), .Y(n572) );
  NOR2XL U1995 ( .A(n1717), .B(n597), .Y(n573) );
  AOI22XL U1996 ( .A0(n57), .A1(n252), .B0(N754), .B1(n253), .Y(n575) );
  AOI211XL U1997 ( .A0(n707), .A1(n652), .B0(n651), .C0(n650), .Y(n653) );
  NOR2XL U1998 ( .A(n659), .B(n703), .Y(n651) );
  NAND2XL U1999 ( .A(n776), .B(write_addr[11]), .Y(n338) );
  AOI211XL U2000 ( .A0(n1364), .A1(n1363), .B0(n1379), .C0(n1398), .Y(n1365)
         );
  XOR2XL U2001 ( .A(\intadd_3/A[7] ), .B(\intadd_3/n3 ), .Y(\intadd_3/SUM[7] )
         );
  INVXL U2002 ( .A(n648), .Y(n652) );
  AOI211XL U2003 ( .A0(N634), .A1(n252), .B0(n569), .C0(n568), .Y(n570) );
  NAND2XL U2004 ( .A(N755), .B(n253), .Y(n566) );
  INVXL U2005 ( .A(n1716), .Y(n567) );
  NOR2XL U2006 ( .A(n571), .B(n234), .Y(n569) );
  AOI211XL U2007 ( .A0(n102), .A1(n649), .B0(n646), .C0(n645), .Y(n647) );
  NOR2XL U2008 ( .A(n654), .B(n703), .Y(n646) );
  XOR2XL U2009 ( .A(\intadd_3/A[8] ), .B(n177), .Y(\intadd_3/SUM[8] ) );
  INVXL U2010 ( .A(n1383), .Y(n1376) );
  OAI211XL U2011 ( .A0(n612), .A1(n636), .B0(n565), .C0(n564), .Y(\C169/Z_14 )
         );
  NOR3XL U2012 ( .A(n597), .B(n1717), .C(n1718), .Y(n563) );
  AOI22XL U2013 ( .A0(N635), .A1(n252), .B0(N756), .B1(n253), .Y(n565) );
  AOI211XL U2014 ( .A0(n89), .A1(n649), .B0(n642), .C0(n641), .Y(n643) );
  NOR2XL U2015 ( .A(n648), .B(n703), .Y(n642) );
  NAND2XL U2016 ( .A(n776), .B(n89), .Y(n341) );
  AOI211XL U2017 ( .A0(n1381), .A1(n1380), .B0(n1387), .C0(n1398), .Y(n1382)
         );
  AND2XL U2018 ( .A(\intadd_3/A[8] ), .B(n177), .Y(n179) );
  AND2XL U2019 ( .A(\intadd_3/A[7] ), .B(\intadd_3/n3 ), .Y(n177) );
  INVXL U2020 ( .A(n1300), .Y(\intadd_3/A[1] ) );
  INVXL U2021 ( .A(\intadd_3/SUM[0] ), .Y(n1425) );
  NOR2XL U2022 ( .A(n1415), .B(n1412), .Y(n1292) );
  INVXL U2023 ( .A(n1287), .Y(n1161) );
  NAND2XL U2024 ( .A(n2136), .B(\next_cr_y[0] ), .Y(n1162) );
  INVXL U2025 ( .A(n1160), .Y(n2136) );
  NAND2XL U2026 ( .A(n1283), .B(n1155), .Y(n1291) );
  NAND2XL U2027 ( .A(n1289), .B(\intadd_3/A[0] ), .Y(n1288) );
  AND2XL U2028 ( .A(n1284), .B(\next_cr_y[0] ), .Y(n1294) );
  NAND2XL U2029 ( .A(n1149), .B(n1148), .Y(n1154) );
  INVXL U2030 ( .A(n1143), .Y(n1151) );
  NOR2XL U2031 ( .A(n1297), .B(n2134), .Y(n1136) );
  INVXL U2032 ( .A(n1134), .Y(n1137) );
  INVXL U2033 ( .A(n1129), .Y(n1132) );
  AND3XL U2034 ( .A(n1125), .B(n1124), .C(\intadd_3/A[0] ), .Y(n1127) );
  NAND2XL U2035 ( .A(n1124), .B(\intadd_3/A[0] ), .Y(n1118) );
  NOR2XL U2036 ( .A(n1119), .B(n1305), .Y(n1121) );
  INVXL U2037 ( .A(n1114), .Y(n1117) );
  NAND2XL U2038 ( .A(n1126), .B(n1131), .Y(n1130) );
  NAND3XL U2039 ( .A(n1128), .B(n1125), .C(n1124), .Y(n1126) );
  OAI211XL U2040 ( .A0(n1104), .A1(n1120), .B0(n1103), .C0(n1102), .Y(n1105)
         );
  NAND2XL U2041 ( .A(n1101), .B(n1308), .Y(n1102) );
  NAND2XL U2042 ( .A(n1119), .B(n1305), .Y(n1120) );
  NOR2XL U2043 ( .A(n1101), .B(n1308), .Y(n1104) );
  INVXL U2044 ( .A(n1097), .Y(n1100) );
  NAND2XL U2045 ( .A(n1116), .B(n1111), .Y(n1115) );
  NAND3XL U2046 ( .A(n1110), .B(n1113), .C(n1107), .Y(n1111) );
  INVXL U2047 ( .A(n1109), .Y(n1107) );
  NAND2XL U2048 ( .A(n1091), .B(n1308), .Y(n1106) );
  AND3XL U2049 ( .A(n1096), .B(n1094), .C(n1308), .Y(n1089) );
  INVXL U2050 ( .A(n1058), .Y(n1061) );
  NAND2XL U2051 ( .A(n1099), .B(n1088), .Y(n1098) );
  NAND3XL U2052 ( .A(n1096), .B(n1090), .C(n1094), .Y(n1088) );
  AND3XL U2053 ( .A(n1056), .B(n1054), .C(next_cr_x[5]), .Y(n1049) );
  XOR2XL U2054 ( .A(n248), .B(next_cr_x[6]), .Y(\DP_OP_719J1_125_1438/n26 ) );
  XOR2XL U2055 ( .A(\next_cr_y[0] ), .B(next_cr_x[5]), .Y(n248) );
  MXI2XL U2056 ( .A(n249), .B(n250), .S0(next_cr_x[5]), .Y(
        \DP_OP_719J1_125_1438/n25 ) );
  NAND2BXL U2057 ( .AN(\next_cr_y[0] ), .B(next_cr_x[6]), .Y(n250) );
  NAND2XL U2058 ( .A(next_cr_x[6]), .B(\next_cr_y[0] ), .Y(n249) );
  INVXL U2059 ( .A(n1310), .Y(n1311) );
  AND2XL U2060 ( .A(next_cr_x[5]), .B(\next_cr_y[0] ), .Y(n186) );
  NAND2XL U2061 ( .A(n1284), .B(n1295), .Y(n1293) );
  INVXL U2062 ( .A(n1000), .Y(n1004) );
  NOR2XL U2063 ( .A(n1310), .B(n997), .Y(n998) );
  INVXL U2064 ( .A(n990), .Y(n992) );
  OAI211XL U2065 ( .A0(write_cntr[1]), .A1(write_cntr[0]), .B0(n131), .C0(n974), .Y(n863) );
  NAND2XL U2066 ( .A(n1048), .B(n1060), .Y(n1059) );
  NAND3XL U2067 ( .A(n1050), .B(n1056), .C(n1054), .Y(n1048) );
  NAND2XL U2068 ( .A(n881), .B(n247), .Y(n855) );
  INVXL U2069 ( .A(n1051), .Y(n247) );
  NAND3XL U2070 ( .A(n869), .B(n867), .C(n859), .Y(n860) );
  INVXL U2071 ( .A(n874), .Y(n862) );
  INVXL U2072 ( .A(n1319), .Y(\intadd_3/A[6] ) );
  NAND2XL U2073 ( .A(n983), .B(n984), .Y(n982) );
  INVXL U2074 ( .A(n981), .Y(n983) );
  NOR2XL U2075 ( .A(n987), .B(n988), .Y(n985) );
  NOR2XL U2076 ( .A(n976), .B(n1361), .Y(n979) );
  INVXL U2077 ( .A(n2137), .Y(n976) );
  NAND2XL U2078 ( .A(write_cntr[1]), .B(write_cntr[0]), .Y(n974) );
  NAND2XL U2079 ( .A(n1360), .B(n1359), .Y(n1357) );
  NAND2XL U2080 ( .A(n1356), .B(n1355), .Y(n1358) );
  NAND2XL U2081 ( .A(n1349), .B(n1348), .Y(n1347) );
  INVXL U2082 ( .A(n1354), .Y(n1360) );
  INVXL U2083 ( .A(n1353), .Y(n1351) );
  NAND2XL U2084 ( .A(n1350), .B(n1349), .Y(n1352) );
  NAND3XL U2085 ( .A(n1346), .B(n1343), .C(n1345), .Y(n1344) );
  NAND2XL U2086 ( .A(n130), .B(n1338), .Y(n1337) );
  NOR2XL U2087 ( .A(n1333), .B(n1334), .Y(n1331) );
  AND2XL U2088 ( .A(n1336), .B(n1334), .Y(n1332) );
  NAND2XL U2089 ( .A(n255), .B(n1329), .Y(n1327) );
  AND2XL U2090 ( .A(n1326), .B(n1325), .Y(n1328) );
  NAND3XL U2091 ( .A(n255), .B(n1326), .C(n1325), .Y(n1323) );
  NAND2XL U2092 ( .A(n1325), .B(n1320), .Y(n1326) );
  INVXL U2093 ( .A(n1329), .Y(n1324) );
  NAND2XL U2094 ( .A(n968), .B(n966), .Y(n967) );
  NAND2XL U2095 ( .A(n965), .B(n84), .Y(n966) );
  INVXL U2096 ( .A(n963), .Y(n968) );
  NAND2XL U2097 ( .A(n2134), .B(n1355), .Y(n960) );
  NAND3XL U2098 ( .A(n963), .B(n84), .C(n962), .Y(n956) );
  INVXL U2099 ( .A(n943), .Y(n946) );
  INVXL U2100 ( .A(n962), .Y(n969) );
  NAND2XL U2101 ( .A(n961), .B(n2134), .Y(n962) );
  OAI2BB2XL U2102 ( .B0(n950), .B1(n949), .A0N(n950), .A1N(n949), .Y(n964) );
  NAND3XL U2103 ( .A(n936), .B(n1345), .C(n935), .Y(n934) );
  NOR2XL U2104 ( .A(n945), .B(n955), .Y(n944) );
  INVXL U2105 ( .A(n953), .Y(n945) );
  NAND2XL U2106 ( .A(write_cntr[4]), .B(write_cntr[3]), .Y(n932) );
  NAND2XL U2107 ( .A(write_cntr[3]), .B(n957), .Y(n952) );
  NAND2BXL U2108 ( .AN(n65), .B(n923), .Y(n927) );
  NOR2BXL U2109 ( .AN(n936), .B(n935), .Y(n929) );
  INVXL U2110 ( .A(n938), .Y(n942) );
  NAND2XL U2111 ( .A(n933), .B(n2139), .Y(n938) );
  NAND3XL U2112 ( .A(n922), .B(n919), .C(n2140), .Y(n920) );
  NOR2XL U2113 ( .A(n1101), .B(n130), .Y(n921) );
  NOR2XL U2114 ( .A(n918), .B(n919), .Y(n1340) );
  NAND2XL U2115 ( .A(n916), .B(n917), .Y(n915) );
  INVXL U2116 ( .A(n914), .Y(n917) );
  AOI21XL U2117 ( .A0(n911), .A1(n908), .B0(n910), .Y(n909) );
  NAND2XL U2118 ( .A(n903), .B(n904), .Y(n902) );
  INVXL U2119 ( .A(n901), .Y(n904) );
  NOR2XL U2120 ( .A(n916), .B(n914), .Y(n905) );
  INVXL U2121 ( .A(n896), .Y(n899) );
  INVXL U2122 ( .A(n895), .Y(n900) );
  INVXL U2123 ( .A(n892), .Y(n897) );
  NOR2XL U2124 ( .A(n891), .B(n255), .Y(n893) );
  NOR2XL U2125 ( .A(n890), .B(n892), .Y(n1330) );
  NAND2XL U2126 ( .A(n888), .B(n889), .Y(n887) );
  INVXL U2127 ( .A(n886), .Y(n889) );
  NOR2XL U2128 ( .A(n901), .B(n903), .Y(n890) );
  INVXL U2129 ( .A(n891), .Y(n2141) );
  NOR2XL U2130 ( .A(n881), .B(n1322), .Y(n884) );
  INVXL U2131 ( .A(n877), .Y(n883) );
  NAND3XL U2132 ( .A(n875), .B(n1320), .C(n874), .Y(n873) );
  NOR2XL U2133 ( .A(n888), .B(n886), .Y(n876) );
  INVXL U2134 ( .A(n872), .Y(n879) );
  NOR2XL U2135 ( .A(n1321), .B(n856), .Y(n871) );
  INVXL U2136 ( .A(n882), .Y(n880) );
  NOR2BXL U2137 ( .AN(n875), .B(n874), .Y(n870) );
  NOR3XL U2138 ( .A(n777), .B(n251), .C(n776), .Y(n845) );
  NAND2XL U2139 ( .A(write_cntr[13]), .B(n848), .Y(n844) );
  AND2XL U2140 ( .A(n2143), .B(n869), .Y(n175) );
  NOR2XL U2141 ( .A(n189), .B(n849), .Y(n846) );
  INVXL U2142 ( .A(n864), .Y(n930) );
  INVXL U2143 ( .A(n852), .Y(n853) );
  AOI32XL U2144 ( .A0(write_cntr[7]), .A1(n857), .A2(n907), .B0(write_cntr[8]), 
        .B1(n857), .Y(n858) );
  INVXL U2145 ( .A(n2930), .Y(n2118) );
  NAND3XL U2146 ( .A(write_cntr[5]), .B(write_cntr[4]), .C(write_cntr[3]), .Y(
        n841) );
  NAND4XL U2147 ( .A(write_cntr[5]), .B(write_cntr[4]), .C(write_cntr[3]), .D(
        n957), .Y(n865) );
  NAND2XL U2148 ( .A(n2121), .B(n777), .Y(n2929) );
  NAND2XL U2149 ( .A(n2322), .B(n840), .Y(n284) );
  NAND3XL U2150 ( .A(write_cntr[8]), .B(write_cntr[7]), .C(write_cntr[6]), .Y(
        n854) );
  AOI211XL U2151 ( .A0(N636), .A1(n252), .B0(n560), .C0(n559), .Y(n561) );
  NAND2XL U2152 ( .A(N757), .B(n253), .Y(n557) );
  NOR2XL U2153 ( .A(n556), .B(n154), .Y(n560) );
  INVXL U2154 ( .A(n562), .Y(n556) );
  NOR2BXL U2155 ( .AN(curr_photo_addr[16]), .B(n718), .Y(\C1/Z_16 ) );
  AOI211XL U2156 ( .A0(n88), .A1(n649), .B0(n638), .C0(n637), .Y(n639) );
  NOR2XL U2157 ( .A(n644), .B(n703), .Y(n638) );
  NAND2XL U2158 ( .A(n776), .B(n88), .Y(n344) );
  NAND2XL U2159 ( .A(n777), .B(n1385), .Y(n345) );
  NAND2XL U2160 ( .A(n1406), .B(n1379), .Y(n1383) );
  OAI211XL U2161 ( .A0(n612), .A1(n2944), .B0(n555), .C0(n554), .Y(\C169/Z_16 ) );
  NOR2XL U2162 ( .A(write_addr[17]), .B(n597), .Y(n552) );
  AOI211XL U2163 ( .A0(N637), .A1(n252), .B0(n550), .C0(n549), .Y(n555) );
  NOR4XL U2164 ( .A(n597), .B(write_addr[18]), .C(n558), .D(n154), .Y(n549) );
  INVXL U2165 ( .A(n551), .Y(n558) );
  AND2XL U2166 ( .A(N758), .B(n253), .Y(n550) );
  NOR2BXL U2167 ( .AN(curr_photo_addr[17]), .B(n718), .Y(\C1/Z_17 ) );
  AOI211XL U2168 ( .A0(write_addr[15]), .A1(n649), .B0(n634), .C0(n633), .Y(
        n635) );
  AOI211XL U2169 ( .A0(n1400), .A1(n1399), .B0(n1405), .C0(n1398), .Y(n1401)
         );
  NAND2BXL U2170 ( .AN(n1396), .B(n1397), .Y(n1399) );
  NOR2XL U2171 ( .A(n1400), .B(n1431), .Y(n1402) );
  NOR2XL U2172 ( .A(n640), .B(n703), .Y(n634) );
  INVXL U2173 ( .A(n777), .Y(n1378) );
  AOI211XL U2174 ( .A0(n1391), .A1(n1392), .B0(n1397), .C0(n1398), .Y(n1393)
         );
  NOR2XL U2175 ( .A(n1388), .B(n235), .Y(n1390) );
  AOI211XL U2176 ( .A0(N638), .A1(n252), .B0(n531), .C0(n522), .Y(n532) );
  NAND2XL U2177 ( .A(N759), .B(n253), .Y(n517) );
  NOR2BXL U2178 ( .AN(n624), .B(n612), .Y(n531) );
  AOI211XL U2179 ( .A0(n769), .A1(n516), .B0(n553), .C0(n515), .Y(n544) );
  INVXL U2180 ( .A(n598), .Y(n515) );
  AOI211XL U2181 ( .A0(n1695), .A1(n1694), .B0(n1693), .C0(n1692), .Y(n1696)
         );
  AOI211XL U2182 ( .A0(n1703), .A1(n1691), .B0(n171), .C0(n1721), .Y(n1693) );
  NAND2XL U2183 ( .A(n772), .B(n207), .Y(n1691) );
  INVXL U2184 ( .A(n623), .Y(n514) );
  NOR2XL U2185 ( .A(read_cntr[0]), .B(n1704), .Y(n1705) );
  INVXL U2186 ( .A(n771), .Y(n1702) );
  NAND2XL U2187 ( .A(n1706), .B(n1699), .Y(n1703) );
  NAND3XL U2188 ( .A(n772), .B(n171), .C(n207), .Y(n510) );
  NAND2BXL U2189 ( .AN(n1711), .B(n1868), .Y(n1712) );
  NOR2BXL U2190 ( .AN(curr_photo_addr[18]), .B(n718), .Y(\C1/Z_18 ) );
  AOI211XL U2191 ( .A0(write_addr[16]), .A1(n649), .B0(n630), .C0(n629), .Y(
        n631) );
  INVXL U2192 ( .A(n1867), .Y(n719) );
  NOR2BXL U2193 ( .AN(n1405), .B(n1404), .Y(n1407) );
  INVXL U2194 ( .A(n1403), .Y(n1408) );
  NOR2XL U2195 ( .A(n636), .B(n703), .Y(n630) );
  INVXL U2196 ( .A(n669), .Y(n710) );
  NAND2XL U2197 ( .A(n776), .B(write_addr[16]), .Y(n349) );
  NAND2XL U2198 ( .A(n777), .B(n1395), .Y(n350) );
  NAND2XL U2199 ( .A(n1406), .B(n1397), .Y(n1394) );
  NAND2XL U2200 ( .A(n1387), .B(n1386), .Y(n1391) );
  NAND2XL U2201 ( .A(n102), .B(n1379), .Y(n1380) );
  INVXL U2202 ( .A(n1362), .Y(n1363) );
  OAI211XL U2203 ( .A0(n167), .A1(n1422), .B0(n1430), .C0(n1432), .Y(n1081) );
  NAND4BXL U2204 ( .AN(n1078), .B(n1403), .C(n1400), .D(n1396), .Y(n1082) );
  AOI211XL U2205 ( .A0(n1364), .A1(n1377), .B0(n1381), .C0(n1718), .Y(n1078)
         );
  INVXL U2206 ( .A(n773), .Y(n1718) );
  INVXL U2207 ( .A(n1075), .Y(n1074) );
  NAND2XL U2208 ( .A(n1073), .B(n102), .Y(n1075) );
  INVXL U2209 ( .A(n1366), .Y(n1367) );
  INVXL U2210 ( .A(n2926), .Y(n283) );
  INVX4 U2211 ( .A(n41), .Y(n257) );
  OAI22X1 U2212 ( .A0(n826), .A1(n831), .B0(n825), .B1(n833), .Y(next_state[2]) );
  NOR2X1 U2213 ( .A(n163), .B(n2949), .Y(n825) );
  INVXL U2214 ( .A(n832), .Y(n826) );
  INVXL U2215 ( .A(n279), .Y(n280) );
  INVXL U2216 ( .A(n836), .Y(n278) );
  OAI21X1 U2217 ( .A0(n148), .A1(n815), .B0(n823), .Y(n832) );
  OAI211XL U2218 ( .A0(n789), .A1(n811), .B0(n788), .C0(global_cntr[11]), .Y(
        n812) );
  AOI211XL U2219 ( .A0(n828), .A1(n204), .B0(n839), .C0(n842), .Y(n829) );
  NAND2XL U2220 ( .A(write_cntr[12]), .B(write_cntr[11]), .Y(n842) );
  NAND4XL U2221 ( .A(n823), .B(n822), .C(n821), .D(n820), .Y(n824) );
  NOR4BXL U2222 ( .AN(n819), .B(n788), .C(n787), .D(n789), .Y(n820) );
  XNOR2X1 U2223 ( .A(n269), .B(global_cntr[9]), .Y(n268) );
  AOI21X1 U2224 ( .A0(n141), .A1(n271), .B0(n270), .Y(n787) );
  AOI21X1 U2225 ( .A0(n144), .A1(n272), .B0(n273), .Y(n786) );
  INVXL U2226 ( .A(n272), .Y(n261) );
  INVXL U2227 ( .A(n260), .Y(n262) );
  AOI21X1 U2228 ( .A0(n143), .A1(n259), .B0(n260), .Y(n800) );
  NOR4XL U2229 ( .A(n793), .B(n790), .C(n794), .D(n795), .Y(n821) );
  AOI21X1 U2230 ( .A0(n138), .A1(n263), .B0(n264), .Y(n794) );
  NOR2XL U2231 ( .A(n792), .B(n791), .Y(n822) );
  INVXL U2232 ( .A(n810), .Y(n265) );
  INVXL U2233 ( .A(n277), .Y(n276) );
  NOR2X2 U2234 ( .A(n818), .B(n810), .Y(n816) );
  NAND3X1 U2235 ( .A(n809), .B(global_cntr[14]), .C(global_cntr[9]), .Y(n810)
         );
  NAND2XL U2236 ( .A(n808), .B(n807), .Y(n1872) );
  INVXL U2237 ( .A(n817), .Y(n275) );
  INVXL U2238 ( .A(n273), .Y(n274) );
  NOR2X1 U2239 ( .A(n143), .B(n259), .Y(n260) );
  NOR2X1 U2240 ( .A(n141), .B(n271), .Y(n270) );
  NAND3X1 U2241 ( .A(n269), .B(global_cntr[10]), .C(global_cntr[9]), .Y(n271)
         );
  NOR2X2 U2242 ( .A(n142), .B(n267), .Y(n269) );
  NAND2XL U2243 ( .A(n2486), .B(n1279), .Y(n1277) );
  INVXL U2244 ( .A(n766), .Y(n622) );
  INVXL U2245 ( .A(n509), .Y(\C169/Z_18 ) );
  NAND2BXL U2246 ( .AN(n1868), .B(n772), .Y(n1698) );
  INVXL U2247 ( .A(n516), .Y(n519) );
  NAND3XL U2248 ( .A(n551), .B(write_addr[17]), .C(write_addr[18]), .Y(n518)
         );
  NAND2XL U2249 ( .A(n773), .B(write_addr[16]), .Y(n508) );
  NAND2XL U2250 ( .A(read_cntr[0]), .B(n1713), .Y(n1720) );
  NOR4XL U2251 ( .A(n1708), .B(n772), .C(write_addr[8]), .D(n1701), .Y(n507)
         );
  NAND2XL U2252 ( .A(n778), .B(read_cntr[0]), .Y(n1701) );
  NAND4XL U2253 ( .A(n1713), .B(n773), .C(n1436), .D(n1435), .Y(n1684) );
  NOR4XL U2254 ( .A(write_addr[17]), .B(write_addr[16]), .C(write_addr[18]), 
        .D(n153), .Y(n1435) );
  NOR3XL U2255 ( .A(write_addr[19]), .B(n207), .C(n1715), .Y(n1436) );
  NAND2XL U2256 ( .A(n102), .B(n89), .Y(n1715) );
  INVXL U2257 ( .A(n772), .Y(n1710) );
  INVX6 U2258 ( .A(n2969), .Y(si_sel) );
  NAND2BXL U2259 ( .AN(curr_photo_size[1]), .B(n778), .Y(n2645) );
  NOR2XL U2260 ( .A(n2955), .B(n1865), .Y(n1866) );
  INVXL U2261 ( .A(n1864), .Y(n2958) );
  OAI211XL U2262 ( .A0(n2493), .A1(n1278), .B0(n1275), .C0(n2476), .Y(n1274)
         );
  INVXL U2263 ( .A(n1273), .Y(n1268) );
  NAND3XL U2264 ( .A(n1273), .B(n2954), .C(n1271), .Y(n1272) );
  NAND2XL U2265 ( .A(n2476), .B(n162), .Y(n2954) );
  NOR2XL U2266 ( .A(work_cntr[4]), .B(n1865), .Y(n1243) );
  NOR2XL U2267 ( .A(n1249), .B(n1253), .Y(n1250) );
  INVXL U2268 ( .A(n1252), .Y(n1256) );
  NAND2XL U2269 ( .A(n1239), .B(n1241), .Y(n1238) );
  INVXL U2270 ( .A(n1241), .Y(n1231) );
  AND3XL U2271 ( .A(n1232), .B(n1228), .C(n1234), .Y(n1240) );
  NAND3XL U2272 ( .A(n1229), .B(n1225), .C(n1230), .Y(n1228) );
  NAND3XL U2273 ( .A(n1212), .B(n1215), .C(n1213), .Y(n1225) );
  INVXL U2274 ( .A(n1219), .Y(n1213) );
  INVXL U2275 ( .A(n1210), .Y(n1208) );
  INVXL U2276 ( .A(n1212), .Y(n1221) );
  NOR2XL U2277 ( .A(n2501), .B(n1201), .Y(n1203) );
  NOR3XL U2278 ( .A(n1194), .B(n1197), .C(n1199), .Y(n1195) );
  NAND2XL U2279 ( .A(n1185), .B(n1184), .Y(n1189) );
  NAND2XL U2280 ( .A(n1180), .B(n1179), .Y(n1185) );
  INVXL U2281 ( .A(n1181), .Y(n1179) );
  NOR2XL U2282 ( .A(n1176), .B(n1201), .Y(n1171) );
  AND2XL U2283 ( .A(n1174), .B(n1182), .Y(n1178) );
  NAND2XL U2284 ( .A(n1169), .B(n1173), .Y(n1174) );
  NAND2XL U2285 ( .A(n1960), .B(n1218), .Y(n1170) );
  INVXL U2286 ( .A(n1863), .Y(n1176) );
  INVXL U2287 ( .A(n1200), .Y(n1194) );
  NAND2XL U2288 ( .A(n1254), .B(n1967), .Y(n1186) );
  NOR2XL U2289 ( .A(work_cntr[13]), .B(n1202), .Y(n1187) );
  NOR2XL U2290 ( .A(n2541), .B(n1865), .Y(n1196) );
  NAND2XL U2291 ( .A(n1227), .B(n193), .Y(n1214) );
  NOR2XL U2292 ( .A(n199), .B(n1047), .Y(n1046) );
  INVXL U2293 ( .A(n2120), .Y(n1047) );
  INVXL U2294 ( .A(n2014), .Y(n1175) );
  AND2XL U2295 ( .A(n2508), .B(n152), .Y(n2647) );
  INVXL U2296 ( .A(n2506), .Y(n2505) );
  OAI21X4 U2297 ( .A0(state[2]), .A1(n32), .B0(n833), .Y(en_so) );
  NOR2XL U2298 ( .A(N205), .B(n1858), .Y(n1860) );
  NAND2XL U2299 ( .A(n1859), .B(n1857), .Y(n1861) );
  AOI22XL U2300 ( .A0(n1856), .A1(n1855), .B0(n1854), .B1(n1853), .Y(n1862) );
  NAND2XL U2301 ( .A(N205), .B(n1858), .Y(n1855) );
  NOR2XL U2302 ( .A(n1854), .B(n1850), .Y(n1851) );
  NAND2XL U2303 ( .A(n1850), .B(n1849), .Y(n1852) );
  MXI2XL U2304 ( .A(n1854), .B(n1853), .S0(n1850), .Y(n1856) );
  INVXL U2305 ( .A(n1844), .Y(n1848) );
  NOR2XL U2306 ( .A(N2283), .B(n1844), .Y(n1841) );
  NAND2XL U2307 ( .A(n52), .B(n1845), .Y(n1842) );
  NAND2XL U2308 ( .A(n1837), .B(n1839), .Y(n1845) );
  NAND2BXL U2309 ( .AN(n1836), .B(n1835), .Y(n1839) );
  NAND2XL U2310 ( .A(n1832), .B(n1831), .Y(n1835) );
  NAND2XL U2311 ( .A(n1836), .B(n1830), .Y(n1837) );
  NAND2XL U2312 ( .A(n1834), .B(n162), .Y(n1830) );
  NAND2XL U2313 ( .A(n1828), .B(n1826), .Y(n1827) );
  NOR2XL U2314 ( .A(work_cntr[4]), .B(n1828), .Y(n1825) );
  NAND2XL U2315 ( .A(n51), .B(n1829), .Y(n1831) );
  NAND2BXL U2316 ( .AN(n1820), .B(n1819), .Y(n1823) );
  NAND2XL U2317 ( .A(n1816), .B(n1815), .Y(n1819) );
  NAND2XL U2318 ( .A(n1814), .B(n1820), .Y(n1821) );
  NAND2XL U2319 ( .A(n1812), .B(n1810), .Y(n1811) );
  NAND2XL U2320 ( .A(n1818), .B(n197), .Y(n1814) );
  NOR2XL U2321 ( .A(work_cntr[6]), .B(n1812), .Y(n1809) );
  NAND2XL U2322 ( .A(n1808), .B(n1813), .Y(n1815) );
  NAND2XL U2323 ( .A(n54), .B(n1803), .Y(n1807) );
  NAND2XL U2324 ( .A(n1800), .B(n1799), .Y(n1803) );
  NOR2XL U2325 ( .A(n129), .B(n1793), .Y(n1798) );
  INVXL U2326 ( .A(n1793), .Y(n1802) );
  NAND2XL U2327 ( .A(n1792), .B(n1791), .Y(n1800) );
  NAND2XL U2328 ( .A(n1797), .B(n193), .Y(n1792) );
  NAND2BXL U2329 ( .AN(n1791), .B(n1794), .Y(n1799) );
  NAND2XL U2330 ( .A(n1787), .B(n1786), .Y(n1790) );
  NAND2XL U2331 ( .A(n1785), .B(n1789), .Y(n1784) );
  INVXL U2332 ( .A(n1777), .Y(n1781) );
  NOR2XL U2333 ( .A(work_cntr[9]), .B(n1785), .Y(n1782) );
  INVXL U2334 ( .A(n1778), .Y(n1774) );
  INVXL U2335 ( .A(n1783), .Y(n1786) );
  NOR2XL U2336 ( .A(work_cntr[10]), .B(n1777), .Y(n1773) );
  NAND2XL U2337 ( .A(n55), .B(n1778), .Y(n1776) );
  NAND2XL U2338 ( .A(n1769), .B(n1771), .Y(n1778) );
  NAND2BXL U2339 ( .AN(n1768), .B(n1767), .Y(n1771) );
  NAND2XL U2340 ( .A(n1764), .B(n1763), .Y(n1767) );
  NAND2XL U2341 ( .A(n1768), .B(n1762), .Y(n1769) );
  NAND2XL U2342 ( .A(n1766), .B(n180), .Y(n1762) );
  NAND2XL U2343 ( .A(n1760), .B(n1758), .Y(n1759) );
  NOR2XL U2344 ( .A(work_cntr[12]), .B(n1760), .Y(n1756) );
  NAND2XL U2345 ( .A(n1757), .B(n1761), .Y(n1763) );
  NAND2BXL U2346 ( .AN(n1752), .B(n1751), .Y(n1755) );
  NAND2XL U2347 ( .A(n1748), .B(n1747), .Y(n1751) );
  NAND2XL U2348 ( .A(n1752), .B(n1746), .Y(n1753) );
  NAND2XL U2349 ( .A(n1750), .B(n184), .Y(n1746) );
  NAND2XL U2350 ( .A(n1744), .B(n1742), .Y(n1743) );
  NOR2XL U2351 ( .A(n256), .B(n1744), .Y(n1741) );
  NAND2XL U2352 ( .A(n1740), .B(n1745), .Y(n1747) );
  INVXL U2353 ( .A(n1735), .Y(n1737) );
  NAND2XL U2354 ( .A(n188), .B(n1739), .Y(n1733) );
  NOR2XL U2355 ( .A(work_cntr[16]), .B(n1727), .Y(n1728) );
  NAND2XL U2356 ( .A(n1734), .B(n188), .Y(n1730) );
  AND2XL U2357 ( .A(n1726), .B(work_cntr[18]), .Y(n1725) );
  NAND2XL U2358 ( .A(n181), .B(n1729), .Y(n1726) );
  NAND2XL U2359 ( .A(n2113), .B(n765), .Y(n621) );
  NOR2X1 U2360 ( .A(n2923), .B(curr_photo_size[1]), .Y(n357) );
  NAND2XL U2361 ( .A(n87), .B(n1686), .Y(n1681) );
  NAND2XL U2362 ( .A(n74), .B(n1682), .Y(n1672) );
  NAND4BXL U2363 ( .AN(n1680), .B(n87), .C(n74), .D(n146), .Y(n1675) );
  NAND2XL U2364 ( .A(n1656), .B(n1655), .Y(n1654) );
  INVXL U2365 ( .A(n1664), .Y(n1652) );
  OAI2BB2XL U2366 ( .B0(n165), .B1(n1646), .A0N(n165), .A1N(n1646), .Y(n1688)
         );
  INVXL U2367 ( .A(n1642), .Y(n1645) );
  NAND2XL U2368 ( .A(n1639), .B(n1638), .Y(n1640) );
  NAND2XL U2369 ( .A(n1637), .B(n1636), .Y(n1638) );
  NAND3XL U2370 ( .A(n1670), .B(n1635), .C(n1666), .Y(n1667) );
  NOR4BXL U2371 ( .AN(n1662), .B(N2282), .C(n1665), .D(n1651), .Y(n1635) );
  NAND2BXL U2372 ( .AN(n1660), .B(n87), .Y(n1651) );
  NOR2BXL U2373 ( .AN(n1657), .B(n1658), .Y(n1685) );
  OAI211XL U2374 ( .A0(n1639), .A1(n1609), .B0(n1611), .C0(n1612), .Y(n1610)
         );
  NAND2BXL U2375 ( .AN(n1608), .B(n1631), .Y(n1639) );
  INVXL U2376 ( .A(n1603), .Y(n1614) );
  AOI22XL U2377 ( .A0(n1605), .A1(n1606), .B0(n1602), .B1(n1601), .Y(n1600) );
  INVXL U2378 ( .A(n1597), .Y(n1602) );
  INVXL U2379 ( .A(n1631), .Y(n1620) );
  NAND2XL U2380 ( .A(n1615), .B(n1595), .Y(n1604) );
  NAND2XL U2381 ( .A(n1618), .B(n1617), .Y(n1595) );
  NOR4BXL U2382 ( .AN(n1605), .B(N2284), .C(n1612), .D(n1596), .Y(n1590) );
  NAND2XL U2383 ( .A(n1625), .B(n1621), .Y(n1608) );
  NAND2XL U2384 ( .A(n1579), .B(n1578), .Y(n1576) );
  INVXL U2385 ( .A(n1575), .Y(n1582) );
  NAND2XL U2386 ( .A(n1597), .B(n1629), .Y(n1596) );
  INVXL U2387 ( .A(n1650), .Y(n1607) );
  AND2XL U2388 ( .A(n1586), .B(n1585), .Y(n1588) );
  NAND2XL U2389 ( .A(n1625), .B(n1632), .Y(n1585) );
  NAND2BXL U2390 ( .AN(n1573), .B(n1571), .Y(n1570) );
  NAND2BXL U2391 ( .AN(n1580), .B(n1589), .Y(n1564) );
  INVXL U2392 ( .A(n1554), .Y(n1556) );
  INVXL U2393 ( .A(n1558), .Y(n1577) );
  NAND2XL U2394 ( .A(n1569), .B(n1597), .Y(n1574) );
  INVXL U2395 ( .A(n1546), .Y(n1543) );
  NAND2XL U2396 ( .A(n1553), .B(n1552), .Y(n1586) );
  NOR4XL U2397 ( .A(n1544), .B(n1535), .C(n1545), .D(n1547), .Y(n1536) );
  NAND2BXL U2398 ( .AN(n1587), .B(n1592), .Y(n1547) );
  NAND3XL U2399 ( .A(n1551), .B(n1569), .C(n197), .Y(n1545) );
  AND2XL U2400 ( .A(n1519), .B(n1530), .Y(n1563) );
  INVXL U2401 ( .A(n1509), .Y(n1511) );
  OAI2BB2XL U2402 ( .B0(n1508), .B1(n1507), .A0N(n1508), .A1N(n1507), .Y(n1529) );
  INVXL U2403 ( .A(n1527), .Y(n1505) );
  NOR4BXL U2404 ( .AN(n1526), .B(work_cntr[6]), .C(n1503), .D(n1535), .Y(n1514) );
  NAND2XL U2405 ( .A(n1559), .B(n1562), .Y(n1535) );
  NAND3XL U2406 ( .A(n1501), .B(n1500), .C(n1520), .Y(n1502) );
  NAND2XL U2407 ( .A(n1519), .B(n1531), .Y(n1520) );
  NAND2BXL U2408 ( .AN(n1492), .B(n1491), .Y(n1493) );
  NAND2XL U2409 ( .A(n1509), .B(n67), .Y(n1495) );
  AOI221XL U2410 ( .A0(n256), .A1(n1490), .B0(n1489), .B1(n1490), .C0(n1492), 
        .Y(n1513) );
  INVXL U2411 ( .A(n1486), .Y(n1489) );
  NAND3XL U2412 ( .A(n194), .B(n1508), .C(n1526), .Y(n1496) );
  INVXL U2413 ( .A(n1483), .Y(n1508) );
  NAND2XL U2414 ( .A(n1481), .B(n1480), .Y(n1482) );
  NAND2XL U2415 ( .A(n1479), .B(n1478), .Y(n1480) );
  NAND2XL U2416 ( .A(work_cntr[10]), .B(n1477), .Y(n1481) );
  NAND2XL U2417 ( .A(n1523), .B(n1532), .Y(n1503) );
  NAND2BXL U2418 ( .AN(n1476), .B(n1533), .Y(n1500) );
  INVXL U2419 ( .A(n1504), .Y(n1484) );
  NAND4XL U2420 ( .A(n1465), .B(n1472), .C(n1464), .D(n193), .Y(n1487) );
  NOR2XL U2421 ( .A(n1490), .B(n1497), .Y(n1464) );
  INVXL U2422 ( .A(n1461), .Y(n1462) );
  NAND2XL U2423 ( .A(n1470), .B(n1469), .Y(n1483) );
  OAI211XL U2424 ( .A0(work_cntr[16]), .A1(n1491), .B0(work_cntr[17]), .C0(
        n1451), .Y(n1452) );
  NAND2XL U2425 ( .A(n1960), .B(n1450), .Y(n1451) );
  NAND2XL U2426 ( .A(n1449), .B(n1460), .Y(n1491) );
  NAND2XL U2427 ( .A(n1461), .B(n2548), .Y(n1501) );
  NAND2XL U2428 ( .A(n1455), .B(n1448), .Y(n1457) );
  NAND2XL U2429 ( .A(n1447), .B(n1454), .Y(n1448) );
  INVXL U2430 ( .A(n2332), .Y(n1450) );
  NOR4XL U2431 ( .A(work_cntr[9]), .B(work_cntr[12]), .C(work_cntr[17]), .D(
        n1458), .Y(n1443) );
  INVXL U2432 ( .A(n1459), .Y(n1449) );
  NAND2XL U2433 ( .A(n1439), .B(n1441), .Y(n1442) );
  NOR3XL U2434 ( .A(work_cntr[13]), .B(work_cntr[15]), .C(n256), .Y(n1439) );
  NOR2XL U2435 ( .A(n256), .B(n1471), .Y(n1440) );
  NAND2BXL U2436 ( .AN(n1445), .B(n1960), .Y(n1437) );
  NAND2XL U2437 ( .A(n161), .B(n182), .Y(n1445) );
  OAI22XL U2438 ( .A0(n2125), .A1(n2124), .B0(n2123), .B1(n2122), .Y(n2126) );
  NOR4XL U2439 ( .A(n140), .B(n1872), .C(n813), .D(n176), .Y(n809) );
  NAND4BBXL U2440 ( .AN(global_cntr[3]), .BN(global_cntr[18]), .C(n1870), .D(
        n176), .Y(n1871) );
  NOR4XL U2441 ( .A(global_cntr[4]), .B(global_cntr[5]), .C(global_cntr[9]), 
        .D(global_cntr[14]), .Y(n1870) );
  OAI22XL U2442 ( .A0(n2953), .A1(n360), .B0(n2952), .B1(n243), .Y(
        next_photo[1]) );
  OAI31XL U2443 ( .A0(cr_read_cntr[3]), .A1(n503), .A2(n478), .B0(n505), .Y(
        N92) );
  AOI221XL U2444 ( .A0(n2963), .A1(n2962), .B0(n2961), .B1(n2962), .C0(n2967), 
        .Y(n2964) );
  OAI22XL U2445 ( .A0(n42), .A1(n246), .B0(n2944), .B1(im_wen_n), .Y(n483) );
  OAI21XL U2446 ( .A0(n40), .A1(n711), .B0(n355), .Y(n530) );
  OAI21XL U2447 ( .A0(n40), .A1(n689), .B0(n331), .Y(n527) );
  OAI21XL U2448 ( .A0(n644), .A1(n40), .B0(n346), .Y(n487) );
  OAI21XL U2449 ( .A0(n40), .A1(n636), .B0(n351), .Y(n485) );
  OAI2BB2XL U2450 ( .B0(n40), .B1(n2133), .A0N(n40), .A1N(write_cntr[2]), .Y(
        n547) );
  OAI22XL U2451 ( .A0(n40), .A1(n2142), .B0(n42), .B1(n204), .Y(n537) );
  OAI22XL U2452 ( .A0(n40), .A1(n874), .B0(n42), .B1(n205), .Y(n533) );
  OAI21XL U2453 ( .A0(n167), .A1(n42), .B0(n334), .Y(n526) );
  OAI22XL U2454 ( .A0(n42), .A1(n208), .B0(im_wen_n), .B1(n353), .Y(n482) );
  OAI21XL U2455 ( .A0(n173), .A1(n2945), .B0(n329), .Y(n529) );
  OAI22XL U2456 ( .A0(n40), .A1(n869), .B0(n2945), .B1(n2144), .Y(n535) );
  OAI22XL U2457 ( .A0(n40), .A1(n2132), .B0(n42), .B1(n201), .Y(n548) );
  OAI22XL U2458 ( .A0(n40), .A1(n2143), .B0(n2945), .B1(n189), .Y(n536) );
  OAI22XL U2459 ( .A0(n40), .A1(n867), .B0(n2945), .B1(n202), .Y(n534) );
  OAI21XL U2460 ( .A0(n40), .A1(n2146), .B0(n335), .Y(n525) );
  OAI21XL U2461 ( .A0(n40), .A1(n2147), .B0(n336), .Y(n524) );
  OAI21XL U2462 ( .A0(n40), .A1(n677), .B0(n337), .Y(n523) );
  OAI21XL U2463 ( .A0(n40), .A1(n668), .B0(n328), .Y(n492) );
  OAI21XL U2464 ( .A0(n664), .A1(n40), .B0(n325), .Y(n491) );
  OAI21XL U2465 ( .A0(n654), .A1(n40), .B0(n340), .Y(n489) );
  OAI21XL U2466 ( .A0(n40), .A1(n648), .B0(n343), .Y(n488) );
  OAI22XL U2467 ( .A0(n2971), .A1(n172), .B0(n151), .B1(n709), .Y(n520) );
  AOI2BB1X1 U2468 ( .A0N(global_cntr[2]), .A1N(n798), .B0(n796), .Y(n797) );
  CLKINVX1 U2469 ( .A(n2660), .Y(n2353) );
  OAI22XL U2470 ( .A0(n2111), .A1(n719), .B0(n2112), .B1(n2967), .Y(n720) );
  AOI221XL U2471 ( .A0(n973), .A1(n205), .B0(n844), .B1(n205), .C0(n845), .Y(
        n866) );
  CLKBUFX3 U2472 ( .A(n775), .Y(n251) );
  OR2X1 U2473 ( .A(n836), .B(n1072), .Y(next_state[1]) );
  AO21X1 U2474 ( .A0(n780), .A1(n834), .B0(n778), .Y(n1072) );
  AOI2BB1X1 U2475 ( .A0N(n190), .A1N(next_state[2]), .B0(n835), .Y(n840) );
  NAND2BX1 U2476 ( .AN(n835), .B(n280), .Y(n2322) );
  NOR2X1 U2477 ( .A(n832), .B(n831), .Y(n836) );
  OAI21XL U2478 ( .A0(n185), .A1(n834), .B0(n833), .Y(n837) );
  NAND3X1 U2479 ( .A(write_cntr[14]), .B(n829), .C(write_cntr[13]), .Y(n2121)
         );
  NOR2X1 U2480 ( .A(n780), .B(en_so), .Y(n779) );
  NOR2X1 U2481 ( .A(n816), .B(n268), .Y(n789) );
  OA21XL U2482 ( .A0(global_cntr[12]), .A1(n270), .B0(n259), .Y(n801) );
  OA21XL U2483 ( .A0(global_cntr[3]), .A1(n796), .B0(n263), .Y(n795) );
  OA21XL U2484 ( .A0(global_cntr[7]), .A1(n266), .B0(n267), .Y(n791) );
  NAND2XL U2485 ( .A(global_cntr[18]), .B(global_cntr[17]), .Y(n813) );
  NOR4XL U2486 ( .A(global_cntr[6]), .B(global_cntr[7]), .C(global_cntr[8]), 
        .D(global_cntr[10]), .Y(n807) );
  NOR4XL U2487 ( .A(global_cntr[11]), .B(global_cntr[12]), .C(global_cntr[13]), 
        .D(global_cntr[15]), .Y(n808) );
  AND2X2 U2488 ( .A(n798), .B(global_cntr[2]), .Y(n796) );
  AOI2BB2X1 U2489 ( .B0(n2111), .B1(n1867), .A0N(n2110), .A1N(n2967), .Y(n620)
         );
  CLKBUFX3 U2490 ( .A(work_cntr[14]), .Y(n256) );
  ADDFXL U2491 ( .A(N2283), .B(n2104), .CI(n2103), .CO(n2105), .S(n2117) );
  NOR2X1 U2492 ( .A(n2932), .B(n284), .Y(n775) );
  OA21XL U2493 ( .A0(n150), .A1(n798), .B0(n2321), .Y(n830) );
  NOR2X1 U2494 ( .A(n818), .B(n139), .Y(n266) );
  NOR2X1 U2495 ( .A(curr_photo_size[0]), .B(n2122), .Y(n1867) );
  CLKINVX1 U2496 ( .A(n827), .Y(n282) );
  AOI2BB1X1 U2497 ( .A0N(global_cntr[1]), .A1N(global_cntr[0]), .B0(n798), .Y(
        \next_glb_cntr[1] ) );
  OAI21XL U2498 ( .A0(n417), .A1(n419), .B0(n425), .Y(n418) );
  OA21XL U2499 ( .A0(curr_time[10]), .A1(n440), .B0(n397), .Y(n399) );
  AO22X1 U2500 ( .A0(n472), .A1(n383), .B0(n470), .B1(n46), .Y(n401) );
  OAI22XL U2501 ( .A0(n378), .A1(n377), .B0(n1029), .B1(n376), .Y(n379) );
  OAI21XL U2502 ( .A0(n435), .A1(n434), .B0(n433), .Y(n436) );
  OAI21XL U2503 ( .A0(curr_time[9]), .A1(n434), .B0(n432), .Y(n433) );
  OAI21XL U2504 ( .A0(n440), .A1(n389), .B0(n393), .Y(n390) );
  OAI22XL U2505 ( .A0(n443), .A1(n429), .B0(n428), .B1(n427), .Y(n430) );
  OAI22XL U2506 ( .A0(n452), .A1(n425), .B0(n424), .B1(n423), .Y(n426) );
  AO22X1 U2507 ( .A0(n472), .A1(n445), .B0(n470), .B1(n444), .Y(n450) );
  OA21XL U2508 ( .A0(n442), .A1(n441), .B0(n440), .Y(n457) );
  OR2X1 U2509 ( .A(n465), .B(n806), .Y(n448) );
  AOI2BB2X1 U2510 ( .B0(n440), .B1(n388), .A0N(n442), .A1N(n389), .Y(n393) );
  OAI21XL U2511 ( .A0(n442), .A1(curr_time[10]), .B0(curr_time[9]), .Y(n396)
         );
  AO21X1 U2512 ( .A0(n2128), .A1(n361), .B0(n2129), .Y(n366) );
  OAI22XL U2513 ( .A0(n1070), .A1(n480), .B0(cr_read_cntr[4]), .B1(n479), .Y(
        n481) );
  OAI21XL U2514 ( .A0(n1069), .A1(n479), .B0(n1070), .Y(n477) );
  OAI2BB1X1 U2515 ( .A0N(n254), .A1N(\C168/DATA3_1 ), .B0(n722), .Y(n723) );
  AOI2BB2X1 U2516 ( .B0(n759), .B1(N1668), .A0N(n756), .A1N(n155), .Y(n722) );
  OAI2BB1X1 U2517 ( .A0N(n760), .A1N(\C168/DATA3_2 ), .B0(n724), .Y(n725) );
  AOI2BB2X1 U2518 ( .B0(n759), .B1(N1669), .A0N(n756), .A1N(n150), .Y(n724) );
  OAI2BB1X1 U2519 ( .A0N(n254), .A1N(\C168/DATA3_3 ), .B0(n726), .Y(n727) );
  AOI2BB2X1 U2520 ( .B0(n759), .B1(N1670), .A0N(n756), .A1N(n156), .Y(n726) );
  OAI2BB1X1 U2521 ( .A0N(n760), .A1N(\C168/DATA3_4 ), .B0(n728), .Y(n729) );
  AOI2BB2X1 U2522 ( .B0(n759), .B1(N1671), .A0N(n756), .A1N(n138), .Y(n728) );
  OAI2BB1X1 U2523 ( .A0N(n254), .A1N(\C168/DATA3_5 ), .B0(n730), .Y(n731) );
  AOI2BB2X1 U2524 ( .B0(n759), .B1(N1672), .A0N(n756), .A1N(n157), .Y(n730) );
  OAI2BB1X1 U2525 ( .A0N(n760), .A1N(\C168/DATA3_6 ), .B0(n732), .Y(n733) );
  AOI2BB2X1 U2526 ( .B0(n759), .B1(N1673), .A0N(n756), .A1N(n139), .Y(n732) );
  OAI2BB1X1 U2527 ( .A0N(n254), .A1N(\C168/DATA3_7 ), .B0(n734), .Y(n735) );
  AOI2BB2X1 U2528 ( .B0(n759), .B1(N1674), .A0N(n756), .A1N(n158), .Y(n734) );
  OAI2BB1X1 U2529 ( .A0N(n760), .A1N(\C168/DATA3_8 ), .B0(n736), .Y(n737) );
  AOI2BB2X1 U2530 ( .B0(n759), .B1(N1675), .A0N(n756), .A1N(n142), .Y(n736) );
  OAI2BB1X1 U2531 ( .A0N(n254), .A1N(\C168/DATA3_9 ), .B0(n738), .Y(n739) );
  AOI2BB2X1 U2532 ( .B0(n759), .B1(N1676), .A0N(n756), .A1N(n147), .Y(n738) );
  OAI2BB1X1 U2533 ( .A0N(n760), .A1N(\C168/DATA3_10 ), .B0(n740), .Y(n741) );
  AOI2BB2X1 U2534 ( .B0(n759), .B1(N1677), .A0N(n756), .A1N(n159), .Y(n740) );
  OAI2BB1X1 U2535 ( .A0N(n254), .A1N(\C168/DATA3_11 ), .B0(n742), .Y(n743) );
  AOI2BB2X1 U2536 ( .B0(n759), .B1(N1678), .A0N(n756), .A1N(n141), .Y(n742) );
  OAI2BB1X1 U2537 ( .A0N(n254), .A1N(\C168/DATA3_12 ), .B0(n744), .Y(n745) );
  AOI2BB2X1 U2538 ( .B0(n759), .B1(N1679), .A0N(n756), .A1N(n174), .Y(n744) );
  OAI2BB1X1 U2539 ( .A0N(n254), .A1N(\C168/DATA3_13 ), .B0(n746), .Y(n747) );
  AOI2BB2X1 U2540 ( .B0(n759), .B1(N1680), .A0N(n756), .A1N(n143), .Y(n746) );
  OAI2BB1X1 U2541 ( .A0N(n254), .A1N(\C168/DATA3_14 ), .B0(n748), .Y(n749) );
  AOI2BB2X1 U2542 ( .B0(n759), .B1(N1681), .A0N(n756), .A1N(n145), .Y(n748) );
  NAND3XL U2543 ( .A(n2638), .B(N2283), .C(n165), .Y(n2636) );
  OAI211XL U2544 ( .A0(n2638), .A1(n165), .B0(n2639), .C0(n199), .Y(n2637) );
  OAI2BB1X1 U2545 ( .A0N(n254), .A1N(\C168/DATA3_15 ), .B0(n750), .Y(n751) );
  AOI2BB2X1 U2546 ( .B0(n759), .B1(N1682), .A0N(n756), .A1N(n144), .Y(n750) );
  OAI2BB1X1 U2547 ( .A0N(n254), .A1N(\C168/DATA3_16 ), .B0(n752), .Y(n753) );
  AOI2BB2X1 U2548 ( .B0(n759), .B1(N1683), .A0N(n756), .A1N(n140), .Y(n752) );
  OAI2BB1X1 U2549 ( .A0N(n254), .A1N(\C168/DATA3_17 ), .B0(n754), .Y(n755) );
  AOI2BB2X1 U2550 ( .B0(n759), .B1(N1684), .A0N(n756), .A1N(n148), .Y(n754) );
  OAI2BB1X1 U2551 ( .A0N(n254), .A1N(\C168/DATA3_18 ), .B0(n757), .Y(n758) );
  AOI2BB2X1 U2552 ( .B0(n759), .B1(N1685), .A0N(n756), .A1N(n149), .Y(n757) );
  OAI22XL U2553 ( .A0(n627), .A1(n103), .B0(n717), .B1(n176), .Y(
        \U3/RSOP_717/C2/Z_19 ) );
  AO22X1 U2554 ( .A0(write_addr[19]), .A1(n628), .B0(n707), .B1(n624), .Y(n625) );
  OAI22XL U2555 ( .A0(n708), .A1(n103), .B0(n717), .B1(n155), .Y(
        \U3/RSOP_717/C2/Z_1 ) );
  OAI22XL U2556 ( .A0(n704), .A1(n212), .B0(n713), .B1(n173), .Y(n705) );
  AO22X1 U2557 ( .A0(curr_photo_addr[1]), .A1(n716), .B0(curr_photo[0]), .B1(
        n780), .Y(n762) );
  AO22X1 U2558 ( .A0(n715), .A1(n714), .B0(n780), .B1(global_cntr[0]), .Y(
        \U3/RSOP_717/C2/Z_0 ) );
  OAI222XL U2559 ( .A0(n212), .A1(n713), .B0(n712), .B1(n711), .C0(n710), .C1(
        n709), .Y(n714) );
  AO22X1 U2560 ( .A0(curr_photo_addr[2]), .A1(n716), .B0(curr_photo[1]), .B1(
        n780), .Y(n763) );
  OAI22XL U2561 ( .A0(n702), .A1(n103), .B0(n717), .B1(n150), .Y(
        \U3/RSOP_717/C2/Z_2 ) );
  OAI22XL U2562 ( .A0(n704), .A1(n173), .B0(n713), .B1(n137), .Y(n699) );
  AO21X1 U2563 ( .A0(curr_photo_addr[3]), .A1(n716), .B0(si_sel), .Y(n764) );
  OAI22XL U2564 ( .A0(n697), .A1(n103), .B0(n717), .B1(n156), .Y(
        \U3/RSOP_717/C2/Z_3 ) );
  OAI22XL U2565 ( .A0(n704), .A1(n137), .B0(n713), .B1(n211), .Y(n694) );
  AO21X1 U2566 ( .A0(curr_photo_addr[4]), .A1(n716), .B0(si_sel), .Y(\C1/Z_4 )
         );
  OAI22XL U2567 ( .A0(n693), .A1(n103), .B0(n717), .B1(n138), .Y(
        \U3/RSOP_717/C2/Z_4 ) );
  OAI22XL U2568 ( .A0(n704), .A1(n211), .B0(n713), .B1(n167), .Y(n690) );
  OAI22XL U2569 ( .A0(n688), .A1(n103), .B0(n717), .B1(n157), .Y(
        \U3/RSOP_717/C2/Z_5 ) );
  OAI22XL U2570 ( .A0(n704), .A1(n167), .B0(n713), .B1(n213), .Y(n686) );
  OAI22XL U2571 ( .A0(n684), .A1(n103), .B0(n717), .B1(n139), .Y(
        \U3/RSOP_717/C2/Z_6 ) );
  OAI22XL U2572 ( .A0(n704), .A1(n213), .B0(n713), .B1(n136), .Y(n681) );
  AO21X1 U2573 ( .A0(curr_photo_addr[7]), .A1(n716), .B0(si_sel), .Y(\C1/Z_7 )
         );
  OAI22XL U2574 ( .A0(n680), .A1(n103), .B0(n717), .B1(n158), .Y(
        \U3/RSOP_717/C2/Z_7 ) );
  OAI22XL U2575 ( .A0(n704), .A1(n136), .B0(n713), .B1(n168), .Y(n678) );
  OAI21XL U2576 ( .A0(write_addr[9]), .A1(n594), .B0(n593), .Y(n595) );
  OAI22XL U2577 ( .A0(n676), .A1(n103), .B0(n717), .B1(n142), .Y(
        \U3/RSOP_717/C2/Z_8 ) );
  OAI22XL U2578 ( .A0(n704), .A1(n168), .B0(n713), .B1(n207), .Y(n673) );
  OAI22XL U2579 ( .A0(n672), .A1(n103), .B0(n717), .B1(n147), .Y(
        \U3/RSOP_717/C2/Z_9 ) );
  AOI222XL U2580 ( .A0(n671), .A1(n707), .B0(n670), .B1(write_addr[9]), .C0(
        n669), .C1(read_cntr[1]), .Y(n672) );
  OAI21XL U2581 ( .A0(n612), .A1(n659), .B0(n588), .Y(\C169/Z_9 ) );
  AO21X1 U2582 ( .A0(N751), .A1(n253), .B0(n585), .Y(n586) );
  OAI22XL U2583 ( .A0(n667), .A1(n103), .B0(n717), .B1(n159), .Y(
        \U3/RSOP_717/C2/Z_10 ) );
  OAI22XL U2584 ( .A0(n704), .A1(n207), .B0(n713), .B1(n169), .Y(n665) );
  AO21X1 U2585 ( .A0(n251), .A1(\intadd_3/SUM[4] ), .B0(n1318), .Y(n675) );
  OAI21XL U2586 ( .A0(n102), .A1(n582), .B0(n581), .Y(n583) );
  AO21X1 U2587 ( .A0(curr_photo_addr[11]), .A1(n716), .B0(si_sel), .Y(
        \C1/Z_11 ) );
  OAI22XL U2588 ( .A0(n663), .A1(n103), .B0(n717), .B1(n141), .Y(
        \U3/RSOP_717/C2/Z_11 ) );
  OAI22XL U2589 ( .A0(n704), .A1(n233), .B0(n713), .B1(n153), .Y(n660) );
  OAI21XL U2590 ( .A0(n1431), .A1(n1370), .B0(n326), .Y(n327) );
  NOR3BXL U2591 ( .AN(n1714), .B(n89), .C(n597), .Y(n576) );
  OAI22XL U2592 ( .A0(n658), .A1(n103), .B0(n717), .B1(n174), .Y(
        \U3/RSOP_717/C2/Z_12 ) );
  OAI22XL U2593 ( .A0(n704), .A1(n169), .B0(n236), .B1(n713), .Y(n655) );
  OAI21XL U2594 ( .A0(n1431), .A1(n1315), .B0(n323), .Y(n324) );
  OAI21XL U2595 ( .A0(n88), .A1(n573), .B0(n572), .Y(n574) );
  AO21X1 U2596 ( .A0(curr_photo_addr[13]), .A1(n716), .B0(si_sel), .Y(
        \C1/Z_13 ) );
  OAI22XL U2597 ( .A0(n653), .A1(n103), .B0(n717), .B1(n143), .Y(
        \U3/RSOP_717/C2/Z_13 ) );
  OAI22XL U2598 ( .A0(n704), .A1(n153), .B0(n713), .B1(n206), .Y(n650) );
  OAI21XL U2599 ( .A0(n1431), .A1(n1364), .B0(n338), .Y(n339) );
  OAI21XL U2600 ( .A0(n612), .A1(n640), .B0(n570), .Y(\C169/Z_13 ) );
  OAI31XL U2601 ( .A0(n597), .A1(write_addr[15]), .A2(n567), .B0(n566), .Y(
        n568) );
  OA21XL U2602 ( .A0(n1716), .A1(n597), .B0(n598), .Y(n571) );
  AO21X1 U2603 ( .A0(curr_photo_addr[14]), .A1(n716), .B0(si_sel), .Y(
        \C1/Z_14 ) );
  OAI22XL U2604 ( .A0(n647), .A1(n103), .B0(n717), .B1(n145), .Y(
        \U3/RSOP_717/C2/Z_14 ) );
  OAI22XL U2605 ( .A0(n644), .A1(n712), .B0(n713), .B1(n235), .Y(n645) );
  OAI21XL U2606 ( .A0(write_addr[16]), .A1(n563), .B0(n562), .Y(n564) );
  AO21X1 U2607 ( .A0(curr_photo_addr[15]), .A1(n716), .B0(si_sel), .Y(
        \C1/Z_15 ) );
  OAI22XL U2608 ( .A0(n643), .A1(n103), .B0(n717), .B1(n144), .Y(
        \U3/RSOP_717/C2/Z_15 ) );
  OAI22XL U2609 ( .A0(n640), .A1(n712), .B0(n713), .B1(n234), .Y(n641) );
  OAI21XL U2610 ( .A0(n1431), .A1(n1381), .B0(n341), .Y(n342) );
  CLKBUFX3 U2611 ( .A(n1330), .Y(n255) );
  OAI21XL U2612 ( .A0(n612), .A1(n632), .B0(n561), .Y(\C169/Z_15 ) );
  OAI31XL U2613 ( .A0(n597), .A1(write_addr[17]), .A2(n558), .B0(n557), .Y(
        n559) );
  OAI22XL U2614 ( .A0(n639), .A1(n103), .B0(n717), .B1(n140), .Y(
        \U3/RSOP_717/C2/Z_16 ) );
  OAI22XL U2615 ( .A0(n636), .A1(n712), .B0(n713), .B1(n239), .Y(n637) );
  OAI31XL U2616 ( .A0(n553), .A1(n552), .A2(n562), .B0(write_addr[18]), .Y(
        n554) );
  OAI22XL U2617 ( .A0(n635), .A1(n103), .B0(n717), .B1(n148), .Y(
        \U3/RSOP_717/C2/Z_17 ) );
  OAI22XL U2618 ( .A0(n632), .A1(n712), .B0(n713), .B1(n154), .Y(n633) );
  AO21X1 U2619 ( .A0(write_addr[17]), .A1(n776), .B0(n1401), .Y(n352) );
  AOI2BB2X1 U2620 ( .B0(n776), .B1(write_addr[15]), .A0N(n1431), .A1N(n1392), 
        .Y(n347) );
  OAI21XL U2621 ( .A0(n544), .A1(n208), .B0(n532), .Y(\C169/Z_17 ) );
  OAI31XL U2622 ( .A0(n597), .A1(n519), .A2(n518), .B0(n517), .Y(n522) );
  OAI2BB1X1 U2623 ( .A0N(n510), .A1N(n1709), .B0(n778), .Y(n511) );
  AOI2BB2X1 U2624 ( .B0(n619), .B1(n1712), .A0N(n623), .A1N(n513), .Y(n512) );
  OR2X1 U2625 ( .A(n778), .B(write_addr[8]), .Y(n513) );
  OAI22XL U2626 ( .A0(n631), .A1(n103), .B0(n717), .B1(n149), .Y(
        \U3/RSOP_717/C2/Z_18 ) );
  OAI2BB2XL U2627 ( .B0(n2944), .B1(n712), .A0N(write_addr[18]), .A1N(n628), 
        .Y(n629) );
  AOI2BB1X1 U2628 ( .A0N(n1079), .A1N(N748), .B0(n1683), .Y(n774) );
  OA21XL U2629 ( .A0(global_cntr[5]), .A1(n264), .B0(n818), .Y(n793) );
  AOI222XL U2630 ( .A0(n252), .A1(N639), .B0(n519), .B1(n769), .C0(n253), .C1(
        N760), .Y(n509) );
  OAI21XL U2631 ( .A0(n1698), .A1(n172), .B0(n1697), .Y(n613) );
  OR2X1 U2632 ( .A(n518), .B(n208), .Y(n516) );
  AO21X1 U2633 ( .A0(read_cntr[1]), .A1(n1711), .B0(n507), .Y(n614) );
  OR2X1 U2634 ( .A(n2931), .B(n2929), .Y(n151) );
  OA21XL U2635 ( .A0(n792), .A1(n791), .B0(n790), .Y(n811) );
  OAI2BB1X1 U2636 ( .A0N(n819), .A1N(n812), .B0(n785), .Y(n815) );
  NOR2X1 U2637 ( .A(n817), .B(n813), .Y(n814) );
  NOR2X1 U2638 ( .A(n783), .B(n782), .Y(n823) );
  OAI31XL U2639 ( .A0(write_cntr[7]), .A1(write_cntr[5]), .A2(write_cntr[6]), 
        .B0(write_cntr[8]), .Y(n828) );
  AOI2BB2X1 U2640 ( .B0(write_cntr[13]), .B1(n848), .A0N(write_cntr[13]), 
        .A1N(n848), .Y(n843) );
  AO22X1 U2641 ( .A0(write_cntr[13]), .A1(n930), .B0(n843), .B1(n131), .Y(n868) );
  OAI21XL U2642 ( .A0(write_cntr[12]), .A1(n846), .B0(n131), .Y(n847) );
  AOI2BB2X1 U2643 ( .B0(n849), .B1(write_cntr[11]), .A0N(n849), .A1N(
        write_cntr[11]), .Y(n850) );
  AOI2BB2X1 U2644 ( .B0(n1320), .B1(n2143), .A0N(n1320), .A1N(n2143), .Y(n885)
         );
  OAI21XL U2645 ( .A0(n880), .A1(n883), .B0(n879), .Y(n878) );
  AOI2BB2X1 U2646 ( .B0(n2142), .B1(n1325), .A0N(n2142), .A1N(n1325), .Y(n894)
         );
  AOI2BB2X1 U2647 ( .B0(n891), .B1(n255), .A0N(n891), .A1N(n255), .Y(n913) );
  OAI21XL U2648 ( .A0(n900), .A1(n897), .B0(n899), .Y(n898) );
  AOI2BB2X1 U2649 ( .B0(n913), .B1(n912), .A0N(n913), .A1N(n912), .Y(n925) );
  NOR3BXL U2650 ( .AN(n928), .B(n65), .C(n924), .Y(n918) );
  AOI2BB2X1 U2651 ( .B0(n1101), .B1(n130), .A0N(n1101), .A1N(n130), .Y(n933)
         );
  AOI2BB2X1 U2652 ( .B0(n65), .B1(n923), .A0N(n65), .A1N(n923), .Y(n935) );
  OAI21XL U2653 ( .A0(n65), .A1(n924), .B0(n928), .Y(n926) );
  AOI2BB2X1 U2654 ( .B0(n2139), .B1(n1345), .A0N(n2139), .A1N(n1345), .Y(n950)
         );
  AO21X1 U2655 ( .A0(n131), .A1(n931), .B0(n930), .Y(n975) );
  OAI2BB1X1 U2656 ( .A0N(n938), .A1N(n937), .B0(n941), .Y(n939) );
  AOI2BB2X1 U2657 ( .B0(n1350), .B1(n2138), .A0N(n1350), .A1N(n2138), .Y(n961)
         );
  AOI2BB2X1 U2658 ( .B0(n955), .B1(n954), .A0N(n955), .A1N(n953), .Y(n958) );
  OAI21XL U2659 ( .A0(n958), .A1(n1133), .B0(n961), .Y(n959) );
  AOI2BB2X1 U2660 ( .B0(n84), .B1(n965), .A0N(n84), .A1N(n965), .Y(n984) );
  OAI21XL U2661 ( .A0(n972), .A1(n977), .B0(n971), .Y(n970) );
  NAND3BX1 U2662 ( .AN(n977), .B(n980), .C(n2137), .Y(n978) );
  OAI21XL U2663 ( .A0(n1319), .A1(n987), .B0(n988), .Y(n986) );
  OAI21XL U2664 ( .A0(n994), .A1(n1319), .B0(n993), .Y(n991) );
  OAI31XL U2665 ( .A0(n994), .A1(n993), .A2(n992), .B0(n991), .Y(n995) );
  OR2X1 U2666 ( .A(n1006), .B(n1007), .Y(n996) );
  AOI2BB2X1 U2667 ( .B0(n2132), .B1(n1310), .A0N(n2132), .A1N(n1310), .Y(n1163) );
  OA22X1 U2668 ( .A0(n1002), .A1(n1000), .B0(n999), .B1(n998), .Y(n1286) );
  OAI21XL U2669 ( .A0(n1004), .A1(n1310), .B0(n1003), .Y(n1001) );
  OAI21XL U2670 ( .A0(n1310), .A1(n1006), .B0(n1007), .Y(n1005) );
  OR2X1 U2671 ( .A(n1014), .B(curr_time[18]), .Y(n1015) );
  OR2X1 U2672 ( .A(n1030), .B(curr_time[2]), .Y(n1029) );
  NOR2X1 U2673 ( .A(n184), .B(n1037), .Y(n1036) );
  NOR2X1 U2674 ( .A(n188), .B(n1035), .Y(n1034) );
  AO21X1 U2675 ( .A0(n161), .A1(n1031), .B0(n2326), .Y(n2329) );
  OAI2BB1X1 U2676 ( .A0N(n1052), .A1N(next_cr_x[5]), .B0(n1051), .Y(n1053) );
  AOI2BB2X1 U2677 ( .B0(n1056), .B1(n1055), .A0N(n1056), .A1N(n1055), .Y(n1090) );
  AOI2BB2X1 U2678 ( .B0(n1065), .B1(cr_read_cntr[5]), .A0N(n1065), .A1N(n1066), 
        .Y(n1069) );
  AOI2BB2X1 U2679 ( .B0(n208), .B1(n1083), .A0N(n208), .A1N(n1083), .Y(n1410)
         );
  AO21X1 U2680 ( .A0(n1077), .A1(n154), .B0(n1076), .Y(n1400) );
  AO21X1 U2681 ( .A0(n1080), .A1(n136), .B0(n1079), .Y(n1432) );
  OAI21XL U2682 ( .A0(write_addr[8]), .A1(n1084), .B0(n1157), .Y(n1086) );
  AOI2BB2X1 U2683 ( .B0(n1096), .B1(n1095), .A0N(n1096), .A1N(n1095), .Y(n1113) );
  AOI2BB2X1 U2684 ( .B0(n1110), .B1(n1108), .A0N(n1110), .A1N(n1108), .Y(n1128) );
  NOR3BXL U2685 ( .AN(n1110), .B(n1109), .C(n1304), .Y(n1112) );
  AOI2BB2X1 U2686 ( .B0(n1125), .B1(n1118), .A0N(n1125), .A1N(n1118), .Y(n1149) );
  AOI2BB2X1 U2687 ( .B0(n1123), .B1(n1122), .A0N(n1123), .A1N(n1122), .Y(n1146) );
  OAI22XL U2688 ( .A0(n1133), .A1(n1299), .B0(n2134), .B1(n1297), .Y(n1141) );
  AOI2BB2X1 U2689 ( .B0(n1139), .B1(n1138), .A0N(n1139), .A1N(n1138), .Y(n1140) );
  OAI22XL U2690 ( .A0(n1146), .A1(n1147), .B0(n1151), .B1(n1144), .Y(n1145) );
  OAI2BB1X1 U2691 ( .A0N(n1147), .A1N(n1146), .B0(n1145), .Y(n1148) );
  OAI2BB1X1 U2692 ( .A0N(n1152), .A1N(n1151), .B0(n1150), .Y(n1153) );
  AOI2BB2X1 U2693 ( .B0(n1160), .B1(\next_cr_y[0] ), .A0N(n1160), .A1N(
        \next_cr_y[0] ), .Y(n1155) );
  OAI21XL U2694 ( .A0(n1157), .A1(n1398), .B0(n1156), .Y(n1158) );
  AOI2BB2X1 U2695 ( .B0(n1163), .B1(n1162), .A0N(n1285), .A1N(n1161), .Y(n1290) );
  OAI22XL U2696 ( .A0(N742), .A1(n1434), .B0(n173), .B1(n776), .Y(n1164) );
  AO21X1 U2697 ( .A0(n1170), .A1(work_cntr[17]), .B0(n1166), .Y(n1173) );
  AO21X1 U2698 ( .A0(n1962), .A1(n1254), .B0(n152), .Y(n1167) );
  AO21X1 U2699 ( .A0(n1173), .A1(n1172), .B0(n1169), .Y(n1182) );
  OAI222XL U2700 ( .A0(n1180), .A1(n1193), .B0(n1180), .B1(n181), .C0(n1193), 
        .C1(n1179), .Y(n1177) );
  AOI2BB2X1 U2701 ( .B0(n1192), .B1(n1193), .A0N(n1192), .A1N(n1193), .Y(n1191) );
  OAI21XL U2702 ( .A0(n1183), .A1(n1182), .B0(n1181), .Y(n1184) );
  OAI21XL U2703 ( .A0(work_cntr[15]), .A1(n1200), .B0(n1192), .Y(n1188) );
  OAI2BB1X1 U2704 ( .A0N(n2502), .A1N(n1206), .B0(n1199), .Y(n1190) );
  AOI2BB2X1 U2705 ( .B0(n1191), .B1(n1190), .A0N(n1191), .A1N(n1194), .Y(n1204) );
  OAI21XL U2706 ( .A0(n1197), .A1(n1199), .B0(n1200), .Y(n1198) );
  OAI21XL U2707 ( .A0(work_cntr[13]), .A1(n1216), .B0(n1204), .Y(n1205) );
  AO21X1 U2708 ( .A0(n2548), .A1(n1221), .B0(n1217), .Y(n1209) );
  NAND3BX1 U2709 ( .AN(n1211), .B(n1216), .C(n1217), .Y(n1215) );
  AO21X1 U2710 ( .A0(work_cntr[9]), .A1(n1214), .B0(n1218), .Y(n1232) );
  OA21XL U2711 ( .A0(n1217), .A1(n1216), .B0(n1215), .Y(n1222) );
  OAI21XL U2712 ( .A0(work_cntr[11]), .A1(n1229), .B0(n1219), .Y(n1220) );
  AOI2BB1X1 U2713 ( .A0N(work_cntr[10]), .A1N(n1232), .B0(n1230), .Y(n1223) );
  AOI2BB1X1 U2714 ( .A0N(n1234), .A1N(n1232), .B0(n1240), .Y(n1237) );
  OA21XL U2715 ( .A0(n1230), .A1(n1229), .B0(n1228), .Y(n1233) );
  OAI21XL U2716 ( .A0(n1231), .A1(n1232), .B0(n1233), .Y(n1235) );
  OAI21XL U2717 ( .A0(work_cntr[8]), .A1(n1246), .B0(n1239), .Y(n1236) );
  AOI2BB2X1 U2718 ( .B0(n1237), .B1(n1236), .A0N(n1237), .A1N(n1241), .Y(n1244) );
  AOI2BB2X1 U2719 ( .B0(n1247), .B1(n1246), .A0N(n1247), .A1N(n1245), .Y(n1257) );
  OAI21XL U2720 ( .A0(work_cntr[6]), .A1(n1251), .B0(n1257), .Y(n1248) );
  AO21X1 U2721 ( .A0(n1258), .A1(n1259), .B0(n1264), .Y(n1263) );
  OAI21XL U2722 ( .A0(work_cntr[5]), .A1(n1267), .B0(n1258), .Y(n1260) );
  AOI2BB2X1 U2723 ( .B0(n1261), .B1(n1260), .A0N(n1261), .A1N(n1259), .Y(n1266) );
  OA21XL U2724 ( .A0(n1266), .A1(n1264), .B0(n1267), .Y(n1262) );
  AOI2BB2X1 U2725 ( .B0(n1263), .B1(n1267), .A0N(n1263), .A1N(n1262), .Y(n1270) );
  OAI21XL U2726 ( .A0(n1264), .A1(n1266), .B0(n1267), .Y(n1265) );
  OAI21XL U2727 ( .A0(n1268), .A1(n1270), .B0(n2470), .Y(n1269) );
  OAI21XL U2728 ( .A0(n2476), .A1(n2470), .B0(n1270), .Y(n1271) );
  AOI2BB2X1 U2729 ( .B0(n1278), .B1(n2476), .A0N(n1278), .A1N(n2476), .Y(n1282) );
  OAI21XL U2730 ( .A0(n1280), .A1(n1279), .B0(n2493), .Y(n1281) );
  AOI2BB2X1 U2731 ( .B0(n1282), .B1(n2486), .A0N(n1282), .A1N(n1281), .Y(n2963) );
  ADDFXL U2732 ( .A(n1297), .B(n1415), .CI(n1288), .CO(n1427), .S(n1420) );
  OAI2BB2XL U2733 ( .B0(n1411), .B1(n1292), .A0N(n1415), .A1N(n1412), .Y(n1419) );
  AO21X1 U2734 ( .A0(n1304), .A1(n1296), .B0(\intadd_3/B[0] ), .Y(n1418) );
  AOI2BB1X1 U2735 ( .A0N(n1299), .A1N(n1308), .B0(n1303), .Y(\intadd_3/CI ) );
  AOI2BB1X1 U2736 ( .A0N(\intadd_3/A[0] ), .A1N(next_cr_x[5]), .B0(n1307), .Y(
        n1302) );
  ADDFXL U2737 ( .A(n1305), .B(n1303), .CI(n1302), .CO(\intadd_3/A[2] ), .S(
        \intadd_3/B[1] ) );
  AOI2BB1X1 U2738 ( .A0N(n1305), .A1N(next_cr_x[6]), .B0(n1309), .Y(n1306) );
  ADDFXL U2739 ( .A(n1308), .B(n1307), .CI(n1306), .CO(\intadd_3/A[3] ), .S(
        \intadd_3/B[2] ) );
  ADDFXL U2740 ( .A(next_cr_x[5]), .B(n1309), .CI(n1308), .CO(\intadd_3/B[4] ), 
        .S(\intadd_3/B[3] ) );
  ADDFXL U2741 ( .A(n186), .B(next_cr_x[6]), .CI(n1311), .CO(\intadd_3/B[6] ), 
        .S(\intadd_3/B[5] ) );
  OR2X1 U2742 ( .A(n1338), .B(n130), .Y(n1339) );
  AOI2BB2X1 U2743 ( .B0(n1372), .B1(n1373), .A0N(n1372), .A1N(n1361), .Y(
        \intadd_3/A[7] ) );
  AOI2BB2X1 U2744 ( .B0(n1386), .B1(n47), .A0N(n1386), .A1N(n47), .Y(n1385) );
  AOI2BB2X1 U2745 ( .B0(n1396), .B1(n1394), .A0N(n1396), .A1N(n1394), .Y(n1395) );
  AOI2BB2X1 U2746 ( .B0(n1412), .B1(n1411), .A0N(n1412), .A1N(n1411), .Y(n1414) );
  ADDFXL U2747 ( .A(n1420), .B(n1419), .CI(n1418), .CO(n1426), .S(n1421) );
  ADDFXL U2748 ( .A(n1427), .B(n1426), .CI(n1425), .CO(n1300), .S(n1429) );
  AOI2BB2X1 U2749 ( .B0(n251), .B1(\intadd_3/SUM[1] ), .A0N(n1430), .A1N(n1431), .Y(n2146) );
  AOI2BB2X1 U2750 ( .B0(n251), .B1(\intadd_3/SUM[2] ), .A0N(n1432), .A1N(n1431), .Y(n2147) );
  AOI2BB2X1 U2751 ( .B0(work_cntr[16]), .B1(n1442), .A0N(n1444), .A1N(n2332), 
        .Y(n1456) );
  OR2X1 U2752 ( .A(n1724), .B(n1444), .Y(n1453) );
  OA21XL U2753 ( .A0(n1447), .A1(n1455), .B0(n1454), .Y(n1446) );
  AOI2BB1X1 U2754 ( .A0N(n1454), .A1N(n1447), .B0(n1446), .Y(n1468) );
  OR2X1 U2755 ( .A(n1457), .B(n187), .Y(n1469) );
  AOI2BB2X1 U2756 ( .B0(n1460), .B1(n1459), .A0N(n1460), .A1N(n1459), .Y(n1490) );
  OAI2BB1X1 U2757 ( .A0N(n1470), .A1N(n1504), .B0(n1469), .Y(n1478) );
  AOI2BB2X1 U2758 ( .B0(n2502), .B1(n1471), .A0N(n2502), .A1N(n1471), .Y(n1474) );
  OAI21XL U2759 ( .A0(n1475), .A1(n1486), .B0(n1474), .Y(n1473) );
  NOR3BXL U2760 ( .AN(n1499), .B(n1503), .C(n1557), .Y(n1485) );
  OR2X1 U2761 ( .A(n1496), .B(n1512), .Y(n1498) );
  OAI21XL U2762 ( .A0(n1516), .A1(n1511), .B0(n67), .Y(n1510) );
  AO21X1 U2763 ( .A0(n1517), .A1(n1516), .B0(n1515), .Y(n1539) );
  OAI21XL U2764 ( .A0(n1527), .A1(n1525), .B0(n1526), .Y(n1524) );
  AOI2BB1X1 U2765 ( .A0N(n1542), .A1N(n1541), .B0(n1540), .Y(n1573) );
  OR4X1 U2766 ( .A(n1578), .B(n1547), .C(n1633), .D(work_cntr[4]), .Y(n1565)
         );
  OAI21XL U2767 ( .A0(n1575), .A1(n1556), .B0(n1557), .Y(n1555) );
  OAI21XL U2768 ( .A0(n1563), .A1(n1561), .B0(n1562), .Y(n1560) );
  OAI31XL U2769 ( .A0(n1563), .A1(n1562), .A2(n1561), .B0(n1560), .Y(n1572) );
  OA21XL U2770 ( .A0(n1567), .A1(n1598), .B0(n1566), .Y(n1568) );
  AOI2BB2X1 U2771 ( .B0(n1588), .B1(n1587), .A0N(n1588), .A1N(n1587), .Y(n1621) );
  AOI2BB2X1 U2772 ( .B0(n1592), .B1(n1591), .A0N(n1592), .A1N(n1591), .Y(n1593) );
  AOI2BB2X1 U2773 ( .B0(n1594), .B1(n1593), .A0N(n1594), .A1N(n1593), .Y(n1617) );
  OA21XL U2774 ( .A0(n1599), .A1(n1626), .B0(n1598), .Y(n1601) );
  NAND3BX1 U2775 ( .AN(n1660), .B(n1629), .C(n199), .Y(n1622) );
  OA21XL U2776 ( .A0(n1612), .A1(n1611), .B0(n1610), .Y(n1613) );
  OAI21XL U2777 ( .A0(n1615), .A1(n1617), .B0(n1618), .Y(n1616) );
  OAI21XL U2778 ( .A0(n1633), .A1(n1620), .B0(n1621), .Y(n1619) );
  AOI2BB2X1 U2779 ( .B0(n1636), .B1(n1637), .A0N(n1636), .A1N(n1637), .Y(n1670) );
  OA21XL U2780 ( .A0(n1627), .A1(n1657), .B0(n1626), .Y(n1628) );
  AOI2BB2X1 U2781 ( .B0(n1634), .B1(n1633), .A0N(n1634), .A1N(n1633), .Y(n1666) );
  AOI2BB2X1 U2782 ( .B0(n1650), .B1(n1649), .A0N(n1650), .A1N(n1649), .Y(n1656) );
  AOI2BB2X1 U2783 ( .B0(n1660), .B1(n1659), .A0N(n1660), .A1N(n1659), .Y(n1680) );
  NOR3BXL U2784 ( .AN(n1666), .B(n1665), .C(n1664), .Y(n1669) );
  OAI31XL U2785 ( .A0(n1679), .A1(n1675), .A2(n1678), .B0(n1676), .Y(n1671) );
  AOI2BB2X1 U2786 ( .B0(n1676), .B1(n1675), .A0N(n1676), .A1N(n1674), .Y(n1677) );
  AOI2BB2X1 U2787 ( .B0(n75), .B1(n1682), .A0N(n75), .A1N(n1682), .Y(n2965) );
  OAI31XL U2788 ( .A0(n772), .A1(read_cntr[0]), .A2(write_addr[8]), .B0(n1684), 
        .Y(n1694) );
  AOI2BB2X1 U2789 ( .B0(n1686), .B1(n87), .A0N(n1686), .A1N(n87), .Y(n1690) );
  AOI2BB2X1 U2790 ( .B0(N205), .B1(n1687), .A0N(N205), .A1N(n1687), .Y(n2966)
         );
  AOI222XL U2791 ( .A0(n1700), .A1(n1869), .B0(n1700), .B1(n1698), .C0(n1869), 
        .C1(n1710), .Y(n1692) );
  NAND3BX1 U2792 ( .AN(n1701), .B(n1699), .C(n771), .Y(n1697) );
  AOI222XL U2793 ( .A0(n1708), .A1(n1707), .B0(n1708), .B1(n1706), .C0(n1707), 
        .C1(n1705), .Y(n1709) );
  OAI21XL U2794 ( .A0(n233), .A1(n171), .B0(n769), .Y(n1719) );
  OA21XL U2795 ( .A0(work_cntr[19]), .A1(n182), .B0(n1724), .Y(n1729) );
  AOI2BB2X1 U2796 ( .B0(work_cntr[16]), .B1(n1727), .A0N(work_cntr[16]), .A1N(
        n1727), .Y(n1734) );
  OAI21XL U2797 ( .A0(work_cntr[15]), .A1(n1735), .B0(n1734), .Y(n1732) );
  AOI2BB2X1 U2798 ( .B0(work_cntr[15]), .B1(n1739), .A0N(work_cntr[15]), .A1N(
        n1739), .Y(n1744) );
  OR2X1 U2799 ( .A(n1741), .B(n1740), .Y(n1748) );
  OAI2BB1X1 U2800 ( .A0N(n1748), .A1N(n1745), .B0(n2502), .Y(n1742) );
  OAI2BB1X1 U2801 ( .A0N(n1753), .A1N(n1751), .B0(n184), .Y(n1754) );
  OAI21XL U2802 ( .A0(n1751), .A1(work_cntr[13]), .B0(n1750), .Y(n1749) );
  OR2X1 U2803 ( .A(n1757), .B(n1756), .Y(n1764) );
  OAI2BB1X1 U2804 ( .A0N(n1764), .A1N(n1761), .B0(n2548), .Y(n1758) );
  OA21XL U2805 ( .A0(n2548), .A1(n1763), .B0(n1758), .Y(n1766) );
  OAI2BB1X1 U2806 ( .A0N(n1769), .A1N(n1767), .B0(n180), .Y(n1770) );
  OAI21XL U2807 ( .A0(n1767), .A1(work_cntr[11]), .B0(n1766), .Y(n1765) );
  OAI21XL U2808 ( .A0(n1778), .A1(work_cntr[10]), .B0(n1781), .Y(n1779) );
  OA21XL U2809 ( .A0(n187), .A1(n1790), .B0(n1789), .Y(n1797) );
  OAI2BB1X1 U2810 ( .A0N(n1800), .A1N(n1794), .B0(n193), .Y(n1796) );
  OAI21XL U2811 ( .A0(n1794), .A1(work_cntr[8]), .B0(n1797), .Y(n1795) );
  OR2X1 U2812 ( .A(n1798), .B(n54), .Y(n1805) );
  OAI2BB1X1 U2813 ( .A0N(n1805), .A1N(n1803), .B0(n194), .Y(n1806) );
  OAI21XL U2814 ( .A0(n1803), .A1(n129), .B0(n1802), .Y(n1801) );
  OR2X1 U2815 ( .A(n1809), .B(n1808), .Y(n1816) );
  OAI2BB1X1 U2816 ( .A0N(n1816), .A1N(n1813), .B0(n2600), .Y(n1810) );
  OA21XL U2817 ( .A0(n2600), .A1(n1815), .B0(n1810), .Y(n1818) );
  OAI2BB1X1 U2818 ( .A0N(n1821), .A1N(n1819), .B0(n197), .Y(n1822) );
  OAI21XL U2819 ( .A0(n1819), .A1(work_cntr[5]), .B0(n1818), .Y(n1817) );
  OR2X1 U2820 ( .A(n1825), .B(n51), .Y(n1832) );
  OAI2BB1X1 U2821 ( .A0N(n1832), .A1N(n1829), .B0(n164), .Y(n1826) );
  OA21XL U2822 ( .A0(n164), .A1(n1831), .B0(n1826), .Y(n1834) );
  OAI2BB1X1 U2823 ( .A0N(n1837), .A1N(n1835), .B0(n162), .Y(n1838) );
  OAI21XL U2824 ( .A0(n1835), .A1(N2284), .B0(n1834), .Y(n1833) );
  OR2X1 U2825 ( .A(n1841), .B(n52), .Y(n1843) );
  OAI2BB1X1 U2826 ( .A0N(n1843), .A1N(n1845), .B0(n199), .Y(n1847) );
  OAI21XL U2827 ( .A0(n1845), .A1(N2283), .B0(n1848), .Y(n1846) );
  NAND3BX1 U2828 ( .AN(n1887), .B(n1880), .C(n1882), .Y(n1888) );
  OA21XL U2829 ( .A0(n1884), .A1(n1892), .B0(n1883), .Y(n1885) );
  AOI2BB2X1 U2830 ( .B0(n1887), .B1(n1886), .A0N(n1887), .A1N(n1886), .Y(n1900) );
  NAND3BX1 U2831 ( .AN(n1898), .B(n1900), .C(n1896), .Y(n1903) );
  AOI2BB2X1 U2832 ( .B0(n1891), .B1(n1890), .A0N(n1891), .A1N(n1889), .Y(n1901) );
  OA21XL U2833 ( .A0(n1893), .A1(n1908), .B0(n1892), .Y(n1894) );
  AOI2BB2X1 U2834 ( .B0(n1898), .B1(n1897), .A0N(n1898), .A1N(n1897), .Y(n1917) );
  NAND3BX1 U2835 ( .AN(n1913), .B(n1917), .C(n1907), .Y(n1914) );
  OA22X1 U2836 ( .A0(n1904), .A1(n1903), .B0(n1902), .B1(n1901), .Y(n1915) );
  OR2X1 U2837 ( .A(n1949), .B(write_cntr[6]), .Y(n1922) );
  NAND3BX1 U2838 ( .AN(n1921), .B(n1918), .C(n1931), .Y(n1927) );
  AOI2BB2X1 U2839 ( .B0(n1921), .B1(n1920), .A0N(n1919), .A1N(n1927), .Y(n1948) );
  OAI2BB1X1 U2840 ( .A0N(n1924), .A1N(n1923), .B0(n1922), .Y(n1925) );
  AOI2BB2X1 U2841 ( .B0(n1926), .B1(n1925), .A0N(n1926), .A1N(n1925), .Y(n1945) );
  AOI2BB2X1 U2842 ( .B0(n1931), .B1(n1930), .A0N(n1931), .A1N(n1930), .Y(n1943) );
  OAI21XL U2843 ( .A0(n768), .A1(n166), .B0(n1936), .Y(n1937) );
  OA21XL U2844 ( .A0(n1945), .A1(n1946), .B0(n1942), .Y(n1944) );
  OAI2BB1X1 U2845 ( .A0N(n1966), .A1N(work_cntr[16]), .B0(n1961), .Y(n1973) );
  OA21XL U2846 ( .A0(n1979), .A1(n1973), .B0(n1982), .Y(n1965) );
  AO21X1 U2847 ( .A0(work_cntr[18]), .A1(n1963), .B0(n1962), .Y(n1974) );
  OAI21XL U2848 ( .A0(n1965), .A1(n1968), .B0(n1964), .Y(n1972) );
  OAI21XL U2849 ( .A0(n1979), .A1(n1973), .B0(n1982), .Y(n1969) );
  OAI2BB1X1 U2850 ( .A0N(n1978), .A1N(n1977), .B0(n1984), .Y(n1992) );
  OR2X1 U2851 ( .A(n1992), .B(n1991), .Y(n1983) );
  OAI2BB2XL U2852 ( .B0(n1992), .B1(n1991), .A0N(n1992), .A1N(n1991), .Y(n1994) );
  AOI2BB1X1 U2853 ( .A0N(n1996), .A1N(n2548), .B0(n1995), .Y(n2009) );
  OAI21XL U2854 ( .A0(n2012), .A1(n2018), .B0(n2011), .Y(n2013) );
  OAI21XL U2855 ( .A0(n2039), .A1(n2029), .B0(n2031), .Y(n2030) );
  AOI2BB2X1 U2856 ( .B0(n2041), .B1(n2040), .A0N(n2041), .A1N(n2040), .Y(n2049) );
  AOI2BB2X1 U2857 ( .B0(n110), .B1(n2036), .A0N(n110), .A1N(n2036), .Y(n2056)
         );
  OAI21XL U2858 ( .A0(n2045), .A1(n2043), .B0(n2044), .Y(n2042) );
  AOI2BB1X1 U2859 ( .A0N(n2049), .A1N(n2053), .B0(n2048), .Y(n2052) );
  AOI2BB2X1 U2860 ( .B0(n2051), .B1(n2052), .A0N(n2051), .A1N(n2052), .Y(n2060) );
  AOI2BB2X1 U2861 ( .B0(n2062), .B1(n2061), .A0N(n2062), .A1N(n2061), .Y(n2064) );
  OAI21XL U2862 ( .A0(n2075), .A1(n2069), .B0(n2072), .Y(n2070) );
  OR2X1 U2863 ( .A(n2075), .B(n2074), .Y(n2080) );
  OAI21XL U2864 ( .A0(n2081), .A1(n2079), .B0(n2080), .Y(n2078) );
  OAI21XL U2865 ( .A0(n2102), .A1(n199), .B0(n2089), .Y(n2086) );
  AOI221XL U2866 ( .A0(n2086), .A1(n73), .B0(n2085), .B1(n2084), .C0(n2083), 
        .Y(n2087) );
  OAI22XL U2867 ( .A0(n73), .A1(n2090), .B0(n72), .B1(n2089), .Y(n2094) );
  OAI21XL U2868 ( .A0(n2629), .A1(n2104), .B0(n2092), .Y(n2093) );
  OA21XL U2869 ( .A0(n2095), .A1(n2094), .B0(n2093), .Y(n2096) );
  AOI2BB2X1 U2870 ( .B0(n2115), .B1(n2955), .A0N(n2108), .A1N(n2493), .Y(n2098) );
  AOI2BB2X1 U2871 ( .B0(n2117), .B1(n2955), .A0N(n2310), .A1N(n2108), .Y(n2100) );
  AOI2BB2X1 U2872 ( .B0(n2106), .B1(n2105), .A0N(n2106), .A1N(n2105), .Y(n2116) );
  AOI2BB2X1 U2873 ( .B0(n2107), .B1(n162), .A0N(n2107), .A1N(n162), .Y(n2309)
         );
  AOI2BB2X1 U2874 ( .B0(n2116), .B1(n2955), .A0N(n2108), .A1N(n2309), .Y(n2109) );
  OAI22XL U2875 ( .A0(n40), .A1(n2134), .B0(n2945), .B1(n166), .Y(n546) );
  OAI22XL U2876 ( .A0(n40), .A1(n2135), .B0(n42), .B1(n195), .Y(n545) );
  OAI22XL U2877 ( .A0(n40), .A1(n2136), .B0(n2945), .B1(n203), .Y(n543) );
  OAI22XL U2878 ( .A0(n40), .A1(n2137), .B0(n2945), .B1(n200), .Y(n542) );
  OAI22XL U2879 ( .A0(n40), .A1(n2138), .B0(n42), .B1(n198), .Y(n541) );
  OAI22XL U2880 ( .A0(n40), .A1(n2139), .B0(n2945), .B1(n191), .Y(n540) );
  OAI22XL U2881 ( .A0(n40), .A1(n2140), .B0(n42), .B1(n196), .Y(n539) );
  OAI22XL U2882 ( .A0(n40), .A1(n2141), .B0(n2945), .B1(n192), .Y(n538) );
  AO21X1 U2883 ( .A0(next_work_cntr[17]), .A1(n2158), .B0(n2157), .Y(n2173) );
  AOI2BB2X1 U2884 ( .B0(next_work_cntr[15]), .B1(n2167), .A0N(
        next_work_cntr[15]), .A1N(n2167), .Y(n2169) );
  OAI2BB1X1 U2885 ( .A0N(n2170), .A1N(n2169), .B0(n2172), .Y(n2196) );
  OR2X1 U2886 ( .A(n2178), .B(n2177), .Y(n2180) );
  AO21X1 U2887 ( .A0(n76), .A1(n2183), .B0(n2182), .Y(n2185) );
  OAI31XL U2888 ( .A0(n2186), .A1(n2206), .A2(n2196), .B0(n2185), .Y(n2188) );
  AOI2BB1X1 U2889 ( .A0N(n2200), .A1N(n2188), .B0(n2187), .Y(n2192) );
  OAI21XL U2890 ( .A0(n2198), .A1(n2197), .B0(n2202), .Y(n2199) );
  OAI21XL U2891 ( .A0(n2202), .A1(n2209), .B0(n2201), .Y(n2203) );
  OAI21XL U2892 ( .A0(n2210), .A1(n2208), .B0(n2209), .Y(n2207) );
  OAI31XL U2893 ( .A0(n2210), .A1(n2209), .A2(n2208), .B0(n2207), .Y(n2211) );
  OAI2BB1X1 U2894 ( .A0N(n2218), .A1N(next_work_cntr[10]), .B0(n2217), .Y(
        n2228) );
  OAI21XL U2895 ( .A0(n2225), .A1(n2224), .B0(n2223), .Y(n2226) );
  AOI2BB2X1 U2896 ( .B0(n2690), .B1(n2234), .A0N(n2690), .A1N(n2234), .Y(n2245) );
  AOI2BB2X1 U2897 ( .B0(n2243), .B1(n2242), .A0N(n2243), .A1N(n2242), .Y(n2244) );
  NAND3BX1 U2898 ( .AN(n2259), .B(n2247), .C(n2245), .Y(n2249) );
  AOI2BB1X1 U2899 ( .A0N(n2245), .A1N(n2244), .B0(n2248), .Y(n2261) );
  AOI2BB2X1 U2900 ( .B0(n2247), .B1(n2246), .A0N(n2247), .A1N(n2246), .Y(n2250) );
  OAI22XL U2901 ( .A0(n2269), .A1(n2265), .B0(n2256), .B1(n2261), .Y(n2255) );
  AO21X1 U2902 ( .A0(n2256), .A1(n2261), .B0(n2255), .Y(n2267) );
  AO21X1 U2903 ( .A0(n2259), .A1(n2258), .B0(n2257), .Y(n2260) );
  OAI2BB1X1 U2904 ( .A0N(n2267), .A1N(n2261), .B0(n2260), .Y(n2262) );
  OAI21XL U2905 ( .A0(n2276), .A1(n2274), .B0(n2275), .Y(n2273) );
  AOI2BB2X1 U2906 ( .B0(n2280), .B1(n2279), .A0N(n2280), .A1N(n2279), .Y(n2281) );
  OAI21XL U2907 ( .A0(n2290), .A1(n2287), .B0(n2281), .Y(n2282) );
  OAI21XL U2908 ( .A0(n2291), .A1(n2289), .B0(n2290), .Y(n2288) );
  OAI21XL U2909 ( .A0(n2296), .A1(n2293), .B0(n2292), .Y(n2320) );
  AOI2BB1X1 U2910 ( .A0N(n2303), .A1N(n2302), .B0(n2301), .Y(n2306) );
  OAI31XL U2911 ( .A0(n2307), .A1(n2306), .A2(n2305), .B0(n2304), .Y(n2319) );
  NAND3BX1 U2912 ( .AN(n2330), .B(n2312), .C(n2329), .Y(n2313) );
  OAI31XL U2913 ( .A0(n797), .A1(n2323), .A2(n2950), .B0(n2949), .Y(n2324) );
  AOI2BB2X1 U2914 ( .B0(n2333), .B1(n152), .A0N(n2333), .A1N(n2332), .Y(n2341)
         );
  OAI2BB1X1 U2915 ( .A0N(n2345), .A1N(n2338), .B0(n2336), .Y(n2340) );
  OAI21XL U2916 ( .A0(n2338), .A1(n2337), .B0(n2341), .Y(n2339) );
  OR2X1 U2917 ( .A(n2349), .B(n2343), .Y(n2350) );
  OAI2BB1X1 U2918 ( .A0N(n2350), .A1N(n2348), .B0(n2353), .Y(n2351) );
  OAI21XL U2919 ( .A0(n2348), .A1(n2660), .B0(n2347), .Y(n2346) );
  OR2X1 U2920 ( .A(n2355), .B(n2354), .Y(n2364) );
  OAI2BB1X1 U2921 ( .A0N(n2364), .A1N(n2361), .B0(n2356), .Y(n2357) );
  OA21XL U2922 ( .A0(n2356), .A1(n2363), .B0(n2357), .Y(n2366) );
  OAI2BB1X1 U2923 ( .A0N(n2369), .A1N(n2367), .B0(n2372), .Y(n2370) );
  OAI21XL U2924 ( .A0(n2367), .A1(n2652), .B0(n2366), .Y(n2365) );
  OR2X1 U2925 ( .A(n50), .B(n2373), .Y(n2383) );
  OAI2BB1X1 U2926 ( .A0N(n2383), .A1N(n2380), .B0(n2375), .Y(n2376) );
  OA21XL U2927 ( .A0(n2375), .A1(n2382), .B0(n2376), .Y(n2386) );
  OAI2BB1X1 U2928 ( .A0N(n2389), .A1N(n2387), .B0(n2671), .Y(n2390) );
  OAI21XL U2929 ( .A0(n2387), .A1(n2384), .B0(n2386), .Y(n2385) );
  OR2X1 U2930 ( .A(n49), .B(n2392), .Y(n2401) );
  OAI2BB1X1 U2931 ( .A0N(n2401), .A1N(n2398), .B0(n2394), .Y(n2395) );
  OAI2BB1X1 U2932 ( .A0N(n2407), .A1N(n2405), .B0(n2410), .Y(n2408) );
  OAI21XL U2933 ( .A0(n2405), .A1(n2402), .B0(n2404), .Y(n2403) );
  OR2X1 U2934 ( .A(n2412), .B(n2411), .Y(n2421) );
  OAI2BB1X1 U2935 ( .A0N(n2421), .A1N(n2418), .B0(n2413), .Y(n2414) );
  OA21XL U2936 ( .A0(n2413), .A1(n2420), .B0(n2414), .Y(n2424) );
  OAI2BB1X1 U2937 ( .A0N(n2427), .A1N(n2425), .B0(n2430), .Y(n2428) );
  OAI21XL U2938 ( .A0(n2425), .A1(n2422), .B0(n2424), .Y(n2423) );
  OR2X1 U2939 ( .A(n2432), .B(n53), .Y(n2441) );
  OAI2BB1X1 U2940 ( .A0N(n2441), .A1N(n2438), .B0(n2433), .Y(n2434) );
  OAI2BB1X1 U2941 ( .A0N(n2447), .A1N(n2445), .B0(n2450), .Y(n2448) );
  OAI21XL U2942 ( .A0(n2445), .A1(n2442), .B0(n45), .Y(n2443) );
  OR2X1 U2943 ( .A(n2452), .B(n2451), .Y(n2461) );
  OAI2BB1X1 U2944 ( .A0N(n2461), .A1N(n2458), .B0(n2453), .Y(n2454) );
  OAI31XL U2945 ( .A0(n2458), .A1(n2457), .A2(n2456), .B0(n2455), .Y(n2466) );
  OAI2BB1X1 U2946 ( .A0N(n2467), .A1N(n2465), .B0(n2470), .Y(n2468) );
  OAI21XL U2947 ( .A0(n2465), .A1(n2462), .B0(n44), .Y(n2463) );
  OAI21XL U2948 ( .A0(n2477), .A1(n2476), .B0(n2479), .Y(n2478) );
  OA21XL U2949 ( .A0(n2486), .A1(n2488), .B0(n2490), .Y(n2495) );
  AOI2BB1X1 U2950 ( .A0N(n2495), .A1N(N205), .B0(n2489), .Y(n2498) );
  OAI21XL U2951 ( .A0(N205), .A1(n2497), .B0(n2495), .Y(n2496) );
  OAI21XL U2952 ( .A0(n2498), .A1(n2497), .B0(n2496), .Y(n2924) );
  AO21X1 U2953 ( .A0(work_cntr[15]), .A1(n2504), .B0(n2516), .Y(n2520) );
  AOI2BB2X1 U2954 ( .B0(work_cntr[17]), .B1(n2515), .A0N(work_cntr[17]), .A1N(
        n2515), .Y(n2509) );
  AOI222XL U2955 ( .A0(n2520), .A1(n2523), .B0(n2520), .B1(n2525), .C0(n2523), 
        .C1(work_cntr[16]), .Y(n2518) );
  AOI2BB2X1 U2956 ( .B0(n2519), .B1(n2518), .A0N(n2519), .A1N(n2517), .Y(n2530) );
  OR2X1 U2957 ( .A(n2523), .B(n2525), .Y(n2529) );
  OAI21XL U2958 ( .A0(n2527), .A1(n2526), .B0(n2525), .Y(n2528) );
  OAI21XL U2959 ( .A0(work_cntr[15]), .A1(n2545), .B0(n2530), .Y(n2532) );
  OAI21XL U2960 ( .A0(n256), .A1(n2537), .B0(n2544), .Y(n2534) );
  OR2X1 U2961 ( .A(n2539), .B(n2540), .Y(n2549) );
  AO21X1 U2962 ( .A0(n2540), .A1(n2550), .B0(n2562), .Y(n2554) );
  OAI21XL U2963 ( .A0(n2542), .A1(n2544), .B0(n2545), .Y(n2543) );
  OAI21XL U2964 ( .A0(work_cntr[13]), .A1(n2565), .B0(n2549), .Y(n2551) );
  OAI21XL U2965 ( .A0(work_cntr[12]), .A1(n2555), .B0(n2564), .Y(n2553) );
  OR2X1 U2966 ( .A(n2557), .B(n2558), .Y(n2566) );
  AO21X1 U2967 ( .A0(n2558), .A1(n2567), .B0(n2577), .Y(n2571) );
  AO21X1 U2968 ( .A0(work_cntr[10]), .A1(n2560), .B0(n2559), .Y(n2580) );
  OAI21XL U2969 ( .A0(n2562), .A1(n2564), .B0(n2565), .Y(n2563) );
  OAI21XL U2970 ( .A0(work_cntr[11]), .A1(n2580), .B0(n2566), .Y(n2568) );
  OAI21XL U2971 ( .A0(work_cntr[10]), .A1(n2582), .B0(n2579), .Y(n2570) );
  NOR3BXL U2972 ( .AN(n2580), .B(n2579), .C(n2577), .Y(n2573) );
  NAND3BX1 U2973 ( .AN(n2573), .B(n2574), .C(n2582), .Y(n2590) );
  AOI2BB2X1 U2974 ( .B0(work_cntr[8]), .B1(n2575), .A0N(work_cntr[8]), .A1N(
        n2575), .Y(n2587) );
  OAI21XL U2975 ( .A0(n2577), .A1(n2579), .B0(n2580), .Y(n2578) );
  OAI21XL U2976 ( .A0(work_cntr[9]), .A1(n2594), .B0(n2581), .Y(n2584) );
  OAI21XL U2977 ( .A0(work_cntr[8]), .A1(n2597), .B0(n2589), .Y(n2586) );
  AOI2BB1X1 U2978 ( .A0N(n129), .A1N(n2606), .B0(n2596), .Y(n2598) );
  AO21X1 U2979 ( .A0(n2600), .A1(n2615), .B0(n2607), .Y(n2601) );
  OAI21XL U2980 ( .A0(work_cntr[5]), .A1(n2626), .B0(n2613), .Y(n2611) );
  OAI21XL U2981 ( .A0(work_cntr[4]), .A1(n2635), .B0(n2620), .Y(n2618) );
  OAI21XL U2982 ( .A0(n2619), .A1(n2621), .B0(n2616), .Y(n2617) );
  NAND3BX1 U2983 ( .AN(n2621), .B(n2627), .C(n2626), .Y(n2625) );
  OA21XL U2984 ( .A0(n2627), .A1(n2626), .B0(n2625), .Y(n2634) );
  OAI21XL U2985 ( .A0(n2630), .A1(n2635), .B0(n2634), .Y(n2633) );
  AOI2BB2X1 U2986 ( .B0(N2283), .B1(n2639), .A0N(N2283), .A1N(n2639), .Y(n2640) );
  OAI21XL U2987 ( .A0(N2282), .A1(n2643), .B0(n2642), .Y(n2646) );
  AO21X1 U2988 ( .A0(next_work_cntr[10]), .A1(n2653), .B0(n2678), .Y(n2707) );
  OAI21XL U2989 ( .A0(next_work_cntr[15]), .A1(n2662), .B0(n2661), .Y(n2659)
         );
  OAI21XL U2990 ( .A0(n2665), .A1(n2664), .B0(n2663), .Y(n2667) );
  AO22X1 U2991 ( .A0(n2668), .A1(n2667), .B0(n2695), .B1(n2666), .Y(n2718) );
  OAI21XL U2992 ( .A0(n2675), .A1(n2674), .B0(next_work_cntr[15]), .Y(n2673)
         );
  OAI21XL U2993 ( .A0(n2677), .A1(n2676), .B0(next_work_cntr[13]), .Y(n2681)
         );
  AOI2BB1X1 U2994 ( .A0N(n2695), .A1N(n2694), .B0(n2693), .Y(n2719) );
  AO22X1 U2995 ( .A0(n2719), .A1(n2701), .B0(n2700), .B1(n2699), .Y(n2744) );
  OAI21XL U2996 ( .A0(n2708), .A1(n2706), .B0(n2707), .Y(n2705) );
  OAI21XL U2997 ( .A0(n2722), .A1(n2726), .B0(n2727), .Y(n2721) );
  OAI31XL U2998 ( .A0(n2722), .A1(n2727), .A2(n2726), .B0(n2721), .Y(n2723) );
  OR2X1 U2999 ( .A(n2734), .B(n2733), .Y(n2746) );
  NAND3BX1 U3000 ( .AN(n2756), .B(n2753), .C(n2755), .Y(n2740) );
  OAI21XL U3001 ( .A0(n2737), .A1(n2757), .B0(n48), .Y(n2738) );
  OAI2BB1X1 U3002 ( .A0N(n2747), .A1N(n2774), .B0(n2746), .Y(n2748) );
  OAI21XL U3003 ( .A0(n2762), .A1(n2760), .B0(n2761), .Y(n2759) );
  OAI21XL U3004 ( .A0(n2765), .A1(n2774), .B0(n2764), .Y(n2763) );
  OR2X1 U3005 ( .A(n2772), .B(n2829), .Y(n2801) );
  AOI2BB2X1 U3006 ( .B0(n78), .B1(n2777), .A0N(n78), .A1N(n2777), .Y(n2781) );
  AND4X1 U3007 ( .A(n2795), .B(n2811), .C(n2807), .D(n2788), .Y(n2789) );
  OR2X1 U3008 ( .A(n2859), .B(n2806), .Y(n2828) );
  OR2X1 U3009 ( .A(n2800), .B(n2798), .Y(n2832) );
  OAI21XL U3010 ( .A0(n2797), .A1(n2810), .B0(n2811), .Y(n2796) );
  AOI2BB2X1 U3011 ( .B0(next_work_cntr[4]), .B1(n2805), .A0N(next_work_cntr[4]), .A1N(n2805), .Y(n2853) );
  OR4X1 U3012 ( .A(n2838), .B(n2821), .C(n2860), .D(n2809), .Y(n2839) );
  OR2X1 U3013 ( .A(n2823), .B(n2822), .Y(n2837) );
  NOR3BXL U3014 ( .AN(n2882), .B(next_work_cntr[1]), .C(n2868), .Y(n2866) );
  AOI2BB2X1 U3015 ( .B0(n2836), .B1(n2835), .A0N(n2836), .A1N(n2835), .Y(n2841) );
  OAI31XL U3016 ( .A0(next_work_cntr[2]), .A1(n2867), .A2(n2842), .B0(n2874), 
        .Y(n2847) );
  AOI2BB2X1 U3017 ( .B0(n2853), .B1(n2852), .A0N(n2853), .A1N(n2852), .Y(n2855) );
  AOI2BB2X1 U3018 ( .B0(n2859), .B1(n2858), .A0N(n2859), .A1N(n2858), .Y(n2899) );
  OAI21XL U3019 ( .A0(n2862), .A1(n2864), .B0(n2865), .Y(n2861) );
  OR2X1 U3020 ( .A(n2876), .B(n2877), .Y(n2883) );
  OAI22XL U3021 ( .A0(n2882), .A1(n2883), .B0(n2881), .B1(n2880), .Y(n2879) );
  NAND3BX1 U3022 ( .AN(n2916), .B(n2884), .C(n2908), .Y(n2885) );
  AOI2BB2X1 U3023 ( .B0(n2891), .B1(n2890), .A0N(n2891), .A1N(n2890), .Y(n2904) );
  AO21X1 U3024 ( .A0(n2895), .A1(n2894), .B0(n2893), .Y(n2901) );
  AOI2BB2X1 U3025 ( .B0(next_work_cntr[0]), .B1(n2913), .A0N(next_work_cntr[0]), .A1N(n2913), .Y(n2918) );
  AOI221XL U3026 ( .A0(n2918), .A1(n772), .B0(n2917), .B1(n2916), .C0(n2915), 
        .Y(n2919) );
  OAI21XL U3027 ( .A0(n2920), .A1(n2919), .B0(n765), .Y(n2921) );
  OAI221XL U3028 ( .A0(curr_photo_size[0]), .A1(n2924), .B0(n2923), .B1(n2922), 
        .C0(n2921), .Y(n2925) );
  AOI2BB2X1 U3029 ( .B0(curr_photo[1]), .B1(photo_num[1]), .A0N(curr_photo[1]), 
        .A1N(photo_num[1]), .Y(n2948) );
  AOI2BB2X1 U3030 ( .B0(curr_photo[0]), .B1(photo_num[0]), .A0N(curr_photo[0]), 
        .A1N(photo_num[0]), .Y(n2947) );
endmodule


module DPA ( clk, reset, IM_A, IM_Q, IM_D, IM_WEN, CR_A, CR_Q );
  output [19:0] IM_A;
  input [23:0] IM_Q;
  output [23:0] IM_D;
  output [8:0] CR_A;
  input [12:0] CR_Q;
  input clk, reset;
  output IM_WEN;
  wire   n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, im_d_w_19,
         im_d_w_18, im_d_w_9, im_d_w_8, en_si, en_init_time, en_fb_addr,
         en_photo_num, en_curr_photo_size, en_so, si_sel, init_time_mux_sel,
         \sftr_n[1] , \so_mux_sel[1] , \data_path/si_w[0] ,
         \data_path/si_w[1] , \data_path/si_w[2] , \data_path/si_w[3] ,
         \data_path/si_w[4] , \data_path/si_w[5] , \data_path/si_w[6] ,
         \data_path/si_w[7] , \data_path/si_w[8] , \data_path/si_w[9] ,
         \data_path/si_w[10] , \data_path/si_w[11] , \data_path/si_w[12] ,
         \data_path/si_w[13] , \data_path/si_w[14] , \data_path/si_w[15] ,
         \data_path/si_w[16] , \data_path/si_w[17] , \data_path/si_w[18] ,
         \data_path/si_w[19] , \data_path/si_w[20] , \data_path/si_w[21] ,
         \data_path/si_w[22] , \data_path/si_w[23] , n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n141, n144, n145, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n418, \intadd_0/CI , \intadd_0/SUM[6] ,
         \intadd_0/SUM[5] , \intadd_0/SUM[4] , \intadd_0/SUM[3] ,
         \intadd_0/SUM[2] , \intadd_0/SUM[1] , \intadd_0/SUM[0] ,
         \intadd_0/n7 , \intadd_0/n6 , \intadd_0/n5 , \intadd_0/n4 ,
         \intadd_0/n3 , \intadd_0/n2 , \intadd_0/n1 , \intadd_1/CI ,
         \intadd_1/SUM[6] , \intadd_1/SUM[5] , \intadd_1/SUM[4] ,
         \intadd_1/SUM[3] , \intadd_1/SUM[2] , \intadd_1/SUM[1] ,
         \intadd_1/SUM[0] , \intadd_1/n7 , \intadd_1/n6 , \intadd_1/n5 ,
         \intadd_1/n4 , \intadd_1/n3 , \intadd_1/n2 , \intadd_1/n1 ,
         \intadd_2/CI , \intadd_2/SUM[6] , \intadd_2/SUM[5] ,
         \intadd_2/SUM[4] , \intadd_2/SUM[3] , \intadd_2/SUM[2] ,
         \intadd_2/SUM[1] , \intadd_2/SUM[0] , \intadd_2/n7 , \intadd_2/n6 ,
         \intadd_2/n5 , \intadd_2/n4 , \intadd_2/n3 , \intadd_2/n2 ,
         \intadd_2/n1 , n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n445, n447, n449, n451, n453, n455, n457, n459,
         n461, n463, n465, n466, n467, n468, n469, n470, n471, n473, n475,
         n477, n479, n482, n484, n486, n488, n490, n492, n494, n496, n498,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n755;
  wire   [29:28] im_d_w;
  wire   [23:0] curr_time;
  wire   [19:0] fb_addr;
  wire   [1:0] photo_num;
  wire   [19:0] curr_photo_addr;
  wire   [1:0] curr_photo_size;
  wire   [3:0] expand_sel;
  wire   SYNOPSYS_UNCONNECTED__0;

  CONT ctrl_logic ( .clk(clk), .reset(reset), .im_wen_n(IM_WEN), .cr_a(CR_A), 
        .curr_time(curr_time), .fb_addr(fb_addr), .photo_num(photo_num), 
        .curr_photo_addr(curr_photo_addr), .curr_photo_size(curr_photo_size), 
        .en_si(en_si), .en_init_time(en_init_time), .en_fb_addr(en_fb_addr), 
        .en_photo_num(en_photo_num), .en_curr_photo_addr(n468), 
        .en_curr_photo_size(en_curr_photo_size), .en_so(en_so), .si_sel(si_sel), .init_time_mux_sel(init_time_mux_sel), .sftr_n({\sftr_n[1] , 
        SYNOPSYS_UNCONNECTED__0}), .so_mux_sel({\so_mux_sel[1] , n470}), 
        .expand_sel(expand_sel), .\im_a[19]_BAR (n756), .\im_a[18]_BAR (n757), 
        .\im_a[17]_BAR (n758), .\im_a[16]_BAR (n759), .\im_a[15]_BAR (n760), 
        .\im_a[14]_BAR (n761), .\im_a[13]_BAR (n762), .\im_a[12]_BAR (n763), 
        .\im_a[11]_BAR (n764), .\im_a[10]_BAR (n765), .\im_a[9]_BAR (n766), 
        .\im_a[8]_BAR (n767), .\im_a[7]_BAR (n768), .\im_a[6]_BAR (n769), 
        .\im_a[5]_BAR (n770), .\im_a[4]_BAR (n771), .\im_a[3]_BAR (n772), 
        .\im_a[2]_BAR (n773), .\im_a[1]_BAR (n774), .\im_a[0]_BAR (n775) );
  ADDFXL \intadd_0/U3  ( .A(n777), .B(\data_path/si_w[22] ), .CI(\intadd_0/n3 ), .CO(\intadd_0/n2 ), .S(\intadd_0/SUM[5] ) );
  ADDFXL \intadd_1/U3  ( .A(IM_D[14]), .B(\data_path/si_w[14] ), .CI(
        \intadd_1/n3 ), .CO(\intadd_1/n2 ), .S(\intadd_1/SUM[5] ) );
  ADDFXL \intadd_2/U3  ( .A(IM_D[6]), .B(\data_path/si_w[6] ), .CI(
        \intadd_2/n3 ), .CO(\intadd_2/n2 ), .S(\intadd_2/SUM[5] ) );
  DFFSX1 \data_path/si_reg/q_reg[2]  ( .D(n314), .CK(clk), .SN(n546), .Q(n511), 
        .QN(\data_path/si_w[2] ) );
  DFFSX1 \data_path/si_reg/q_reg[4]  ( .D(n313), .CK(clk), .SN(n546), .Q(n510), 
        .QN(\data_path/si_w[4] ) );
  DFFSX1 \data_path/si_reg/q_reg[1]  ( .D(n315), .CK(clk), .SN(n469), .Q(n505), 
        .QN(\data_path/si_w[1] ) );
  DFFSX1 \data_path/si_reg/q_reg[8]  ( .D(n312), .CK(clk), .SN(n546), .Q(n501), 
        .QN(\data_path/si_w[8] ) );
  DFFSX1 \data_path/init_time_reg/q_reg[1]  ( .D(n145), .CK(clk), .SN(n546), 
        .Q(n650), .QN(curr_time[1]) );
  ADDFXL \intadd_1/U7  ( .A(n784), .B(\data_path/si_w[10] ), .CI(\intadd_1/n7 ), .CO(\intadd_1/n6 ), .S(\intadd_1/SUM[1] ) );
  ADDFXL \intadd_1/U2  ( .A(IM_D[15]), .B(\data_path/si_w[15] ), .CI(
        \intadd_1/n2 ), .CO(\intadd_1/n1 ), .S(\intadd_1/SUM[6] ) );
  ADDFXL \intadd_2/U7  ( .A(IM_D[2]), .B(\data_path/si_w[2] ), .CI(
        \intadd_2/n7 ), .CO(\intadd_2/n6 ), .S(\intadd_2/SUM[1] ) );
  ADDFXL \intadd_2/U2  ( .A(IM_D[7]), .B(\data_path/si_w[7] ), .CI(
        \intadd_2/n2 ), .CO(\intadd_2/n1 ), .S(\intadd_2/SUM[6] ) );
  ADDFXL \intadd_0/U7  ( .A(IM_D[18]), .B(\data_path/si_w[18] ), .CI(
        \intadd_0/n7 ), .CO(\intadd_0/n6 ), .S(\intadd_0/SUM[1] ) );
  ADDFXL \intadd_0/U2  ( .A(n776), .B(\data_path/si_w[23] ), .CI(\intadd_0/n2 ), .CO(\intadd_0/n1 ), .S(\intadd_0/SUM[6] ) );
  ADDFXL \intadd_1/U8  ( .A(n785), .B(\data_path/si_w[9] ), .CI(\intadd_1/CI ), 
        .CO(\intadd_1/n7 ), .S(\intadd_1/SUM[0] ) );
  ADDFXL \intadd_2/U8  ( .A(IM_D[1]), .B(\data_path/si_w[1] ), .CI(
        \intadd_2/CI ), .CO(\intadd_2/n7 ), .S(\intadd_2/SUM[0] ) );
  ADDFXL \intadd_0/U8  ( .A(IM_D[17]), .B(\data_path/si_w[17] ), .CI(
        \intadd_0/CI ), .CO(\intadd_0/n7 ), .S(\intadd_0/SUM[0] ) );
  ADDFXL \intadd_1/U6  ( .A(n783), .B(\data_path/si_w[11] ), .CI(\intadd_1/n6 ), .CO(\intadd_1/n5 ), .S(\intadd_1/SUM[2] ) );
  ADDFXL \intadd_1/U5  ( .A(IM_D[12]), .B(\data_path/si_w[12] ), .CI(
        \intadd_1/n5 ), .CO(\intadd_1/n4 ), .S(\intadd_1/SUM[3] ) );
  ADDFXL \intadd_1/U4  ( .A(IM_D[13]), .B(\data_path/si_w[13] ), .CI(
        \intadd_1/n4 ), .CO(\intadd_1/n3 ), .S(\intadd_1/SUM[4] ) );
  ADDFXL \intadd_2/U6  ( .A(IM_D[3]), .B(\data_path/si_w[3] ), .CI(
        \intadd_2/n6 ), .CO(\intadd_2/n5 ), .S(\intadd_2/SUM[2] ) );
  ADDFXL \intadd_2/U5  ( .A(IM_D[4]), .B(\data_path/si_w[4] ), .CI(
        \intadd_2/n5 ), .CO(\intadd_2/n4 ), .S(\intadd_2/SUM[3] ) );
  ADDFXL \intadd_2/U4  ( .A(IM_D[5]), .B(\data_path/si_w[5] ), .CI(
        \intadd_2/n4 ), .CO(\intadd_2/n3 ), .S(\intadd_2/SUM[4] ) );
  ADDFXL \intadd_0/U6  ( .A(n780), .B(\data_path/si_w[19] ), .CI(\intadd_0/n6 ), .CO(\intadd_0/n5 ), .S(\intadd_0/SUM[2] ) );
  ADDFXL \intadd_0/U5  ( .A(n779), .B(\data_path/si_w[20] ), .CI(\intadd_0/n5 ), .CO(\intadd_0/n4 ), .S(\intadd_0/SUM[3] ) );
  ADDFXL \intadd_0/U4  ( .A(n778), .B(\data_path/si_w[21] ), .CI(\intadd_0/n4 ), .CO(\intadd_0/n3 ), .S(\intadd_0/SUM[4] ) );
  DFFRX2 \data_path/init_time_reg/q_reg[17]  ( .D(n322), .CK(clk), .RN(n469), 
        .Q(curr_time[17]), .QN(n507) );
  DFFSX2 \data_path/init_time_reg/q_reg[2]  ( .D(n144), .CK(clk), .SN(n546), 
        .QN(curr_time[2]) );
  DFFRX2 \data_path/init_time_reg/q_reg[9]  ( .D(n330), .CK(clk), .RN(n546), 
        .Q(curr_time[9]), .QN(n530) );
  DFFRX2 \data_path/init_time_reg/q_reg[12]  ( .D(n327), .CK(clk), .RN(n469), 
        .Q(curr_time[12]), .QN(n520) );
  DFFSX2 \data_path/init_time_reg/q_reg[4]  ( .D(n141), .CK(clk), .SN(n546), 
        .QN(curr_time[4]) );
  DFFRX2 \data_path/init_time_reg/q_reg[10]  ( .D(n329), .CK(clk), .RN(n546), 
        .Q(curr_time[10]), .QN(n506) );
  DFFRX2 \data_path/si_reg/q_reg[16]  ( .D(n418), .CK(clk), .RN(n22), .Q(
        \data_path/si_w[16] ) );
  DFFRX2 \data_path/init_time_reg/q_reg[15]  ( .D(n324), .CK(clk), .RN(n22), 
        .Q(curr_time[15]) );
  DFFRX2 \data_path/init_time_reg/q_reg[14]  ( .D(n325), .CK(clk), .RN(n22), 
        .Q(curr_time[14]) );
  DFFRX2 \data_path/init_time_reg/q_reg[7]  ( .D(n332), .CK(clk), .RN(n22), 
        .Q(curr_time[7]) );
  DFFRX2 \data_path/init_time_reg/q_reg[6]  ( .D(n333), .CK(clk), .RN(n22), 
        .Q(curr_time[6]) );
  DFFRX2 \data_path/init_time_reg/q_reg[20]  ( .D(n319), .CK(clk), .RN(n22), 
        .Q(curr_time[20]) );
  DFFSX2 \data_path/si_reg/q_reg[0]  ( .D(n549), .CK(clk), .SN(n546), .Q(n516), 
        .QN(\data_path/si_w[0] ) );
  DFFRX1 \data_path/si_reg/q_reg[23]  ( .D(n369), .CK(clk), .RN(n546), .Q(
        \data_path/si_w[23] ), .QN(n514) );
  DFFRX1 \data_path/si_reg/q_reg[22]  ( .D(n370), .CK(clk), .RN(n22), .Q(
        \data_path/si_w[22] ), .QN(n513) );
  DFFRX1 \data_path/si_reg/q_reg[21]  ( .D(n371), .CK(clk), .RN(n22), .Q(
        \data_path/si_w[21] ), .QN(n512) );
  DFFRX1 \data_path/si_reg/q_reg[20]  ( .D(n372), .CK(clk), .RN(n22), .Q(
        \data_path/si_w[20] ), .QN(n534) );
  DFFRX1 \data_path/si_reg/q_reg[19]  ( .D(n375), .CK(clk), .RN(n22), .Q(
        \data_path/si_w[19] ), .QN(n528) );
  DFFRX1 \data_path/si_reg/q_reg[18]  ( .D(n378), .CK(clk), .RN(n22), .Q(
        \data_path/si_w[18] ), .QN(n526) );
  DFFRX1 \data_path/si_reg/q_reg[17]  ( .D(n381), .CK(clk), .RN(n22), .Q(
        \data_path/si_w[17] ), .QN(n527) );
  DFFRX1 \data_path/si_reg/q_reg[15]  ( .D(n384), .CK(clk), .RN(n22), .Q(
        \data_path/si_w[15] ), .QN(n525) );
  DFFRX1 \data_path/si_reg/q_reg[14]  ( .D(n387), .CK(clk), .RN(n22), .Q(
        \data_path/si_w[14] ), .QN(n529) );
  DFFRX1 \data_path/si_reg/q_reg[13]  ( .D(n390), .CK(clk), .RN(n22), .Q(
        \data_path/si_w[13] ), .QN(n508) );
  DFFRX1 \data_path/photo_num_reg/q_reg[1]  ( .D(n21), .CK(clk), .RN(n22), .Q(
        photo_num[1]), .QN(n10) );
  DFFRX1 \data_path/si_reg/q_reg[12]  ( .D(n393), .CK(clk), .RN(n22), .Q(
        \data_path/si_w[12] ), .QN(n522) );
  DFFRX1 \data_path/si_reg/q_reg[10]  ( .D(n399), .CK(clk), .RN(n22), .Q(
        \data_path/si_w[10] ), .QN(n500) );
  DFFRX1 \data_path/si_reg/q_reg[9]  ( .D(n402), .CK(clk), .RN(n22), .Q(
        \data_path/si_w[9] ), .QN(n523) );
  DFFRX1 \data_path/si_reg/q_reg[7]  ( .D(n405), .CK(clk), .RN(n22), .Q(
        \data_path/si_w[7] ), .QN(n519) );
  DFFRX1 \data_path/si_reg/q_reg[6]  ( .D(n408), .CK(clk), .RN(n22), .Q(
        \data_path/si_w[6] ), .QN(n524) );
  DFFRX1 \data_path/si_reg/q_reg[5]  ( .D(n411), .CK(clk), .RN(n22), .Q(
        \data_path/si_w[5] ), .QN(n509) );
  DFFRX1 \data_path/si_reg/q_reg[3]  ( .D(n414), .CK(clk), .RN(n22), .Q(
        \data_path/si_w[3] ), .QN(n518) );
  DFFRX1 \data_path/curr_photo_size_reg/q_reg[1]  ( .D(n23), .CK(clk), .RN(n22), .Q(curr_photo_size[1]), .QN(n537) );
  DFFRX1 \data_path/curr_photo_size_reg/q_reg[0]  ( .D(n368), .CK(clk), .RN(
        n22), .Q(curr_photo_size[0]), .QN(n515) );
  DFFRX1 \data_path/init_time_reg/q_reg[16]  ( .D(n323), .CK(clk), .RN(n22), 
        .Q(curr_time[16]), .QN(n503) );
  DFFRX1 \data_path/init_time_reg/q_reg[0]  ( .D(n336), .CK(clk), .RN(n22), 
        .Q(curr_time[0]), .QN(n517) );
  DFFRX1 \data_path/init_time_reg/q_reg[23]  ( .D(n316), .CK(clk), .RN(n22), 
        .Q(curr_time[23]), .QN(n504) );
  DFFRX1 \data_path/init_time_reg/q_reg[22]  ( .D(n317), .CK(clk), .RN(n22), 
        .Q(curr_time[22]), .QN(n532) );
  DFFRX1 \data_path/init_time_reg/q_reg[21]  ( .D(n318), .CK(clk), .RN(n22), 
        .Q(curr_time[21]), .QN(n536) );
  DFFRX1 \data_path/init_time_reg/q_reg[18]  ( .D(n321), .CK(clk), .RN(n22), 
        .Q(curr_time[18]), .QN(n521) );
  DFFRX1 \data_path/init_time_reg/q_reg[13]  ( .D(n326), .CK(clk), .RN(n22), 
        .Q(curr_time[13]), .QN(n535) );
  DFFRX1 \data_path/init_time_reg/q_reg[19]  ( .D(n320), .CK(clk), .RN(n22), 
        .Q(curr_time[19]), .QN(n533) );
  DFFRX1 \data_path/init_time_reg/q_reg[3]  ( .D(n335), .CK(clk), .RN(n22), 
        .Q(curr_time[3]), .QN(n531) );
  DFFRX1 \data_path/init_time_reg/q_reg[11]  ( .D(n328), .CK(clk), .RN(n22), 
        .Q(curr_time[11]), .QN(n502) );
  DFFRX1 \data_path/so_reg/q_reg[25]  ( .D(n341), .CK(clk), .RN(n22), .Q(n778), 
        .QN(n453) );
  DFFRX1 \data_path/so_reg/q_reg[24]  ( .D(n342), .CK(clk), .RN(n22), .Q(n779), 
        .QN(n451) );
  DFFRX1 \data_path/so_reg/q_reg[23]  ( .D(n343), .CK(clk), .RN(n22), .Q(n780), 
        .QN(n449) );
  DFFRX1 \data_path/so_reg/q_reg[13]  ( .D(n353), .CK(clk), .RN(n22), .Q(n783), 
        .QN(n447) );
  DFFRX1 \data_path/so_reg/q_reg[12]  ( .D(n354), .CK(clk), .RN(n22), .Q(n784), 
        .QN(n445) );
  DFFRX1 \data_path/so_reg/q_reg[11]  ( .D(n355), .CK(clk), .RN(n22), .Q(n785), 
        .QN(n443) );
  DFFRX1 \data_path/so_reg/q_reg[28]  ( .D(n338), .CK(clk), .RN(n22), .Q(
        im_d_w[28]), .QN(n539) );
  DFFRX1 \data_path/so_reg/q_reg[18]  ( .D(n348), .CK(clk), .RN(n22), .Q(
        im_d_w_18), .QN(n540) );
  DFFRX1 \data_path/so_reg/q_reg[8]  ( .D(n358), .CK(clk), .RN(n22), .Q(
        im_d_w_8), .QN(n538) );
  DFFRX1 \data_path/so_reg/q_reg[26]  ( .D(n340), .CK(clk), .RN(n22), .Q(n777), 
        .QN(n455) );
  DFFRX1 \data_path/so_reg/q_reg[27]  ( .D(n339), .CK(clk), .RN(n22), .Q(n776), 
        .QN(n457) );
  DFFRX1 \data_path/so_reg/q_reg[20]  ( .D(n346), .CK(clk), .RN(n22), .Q(n782), 
        .QN(n463) );
  DFFRX1 \data_path/so_reg/q_reg[0]  ( .D(n366), .CK(clk), .RN(n22), .Q(n787), 
        .QN(n461) );
  DFFRX1 \data_path/so_reg/q_reg[10]  ( .D(n356), .CK(clk), .RN(n22), .Q(n786), 
        .QN(n459) );
  DFFRX1 \data_path/photo_num_reg/q_reg[0]  ( .D(n367), .CK(clk), .RN(n469), 
        .Q(photo_num[0]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[0]  ( .D(n415), .CK(clk), .RN(
        n546), .Q(curr_photo_addr[0]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[2]  ( .D(n17), .CK(clk), .RN(
        n469), .Q(curr_photo_addr[2]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[15]  ( .D(n382), .CK(clk), .RN(
        n546), .Q(curr_photo_addr[15]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[14]  ( .D(n385), .CK(clk), .RN(
        n469), .Q(curr_photo_addr[14]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[4]  ( .D(n15), .CK(clk), .RN(
        n546), .Q(curr_photo_addr[4]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[19]  ( .D(n373), .CK(clk), .RN(
        n546), .Q(curr_photo_addr[19]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[18]  ( .D(n376), .CK(clk), .RN(
        n469), .Q(curr_photo_addr[18]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[17]  ( .D(n379), .CK(clk), .RN(
        n469), .Q(curr_photo_addr[17]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[9]  ( .D(n400), .CK(clk), .RN(
        n546), .Q(curr_photo_addr[9]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[6]  ( .D(n406), .CK(clk), .RN(
        n469), .Q(curr_photo_addr[6]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[12]  ( .D(n391), .CK(clk), .RN(
        n546), .Q(curr_photo_addr[12]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[10]  ( .D(n397), .CK(clk), .RN(
        n546), .Q(curr_photo_addr[10]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[5]  ( .D(n409), .CK(clk), .RN(
        n469), .Q(curr_photo_addr[5]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[1]  ( .D(n19), .CK(clk), .RN(
        n469), .Q(curr_photo_addr[1]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[8]  ( .D(n13), .CK(clk), .RN(
        n546), .Q(curr_photo_addr[8]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[7]  ( .D(n403), .CK(clk), .RN(
        n546), .Q(curr_photo_addr[7]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[3]  ( .D(n412), .CK(clk), .RN(
        n469), .Q(curr_photo_addr[3]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[13]  ( .D(n388), .CK(clk), .RN(
        n469), .Q(curr_photo_addr[13]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[11]  ( .D(n394), .CK(clk), .RN(
        n546), .Q(curr_photo_addr[11]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[16]  ( .D(n11), .CK(clk), .RN(
        n546), .Q(curr_photo_addr[16]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[16]  ( .D(n12), .CK(clk), .RN(n546), .Q(
        fb_addr[16]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[19]  ( .D(n374), .CK(clk), .RN(n546), 
        .Q(fb_addr[19]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[18]  ( .D(n377), .CK(clk), .RN(n546), 
        .Q(fb_addr[18]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[17]  ( .D(n380), .CK(clk), .RN(n469), 
        .Q(fb_addr[17]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[15]  ( .D(n383), .CK(clk), .RN(n546), 
        .Q(fb_addr[15]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[12]  ( .D(n392), .CK(clk), .RN(n469), 
        .Q(fb_addr[12]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[6]  ( .D(n407), .CK(clk), .RN(n469), .Q(
        fb_addr[6]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[5]  ( .D(n410), .CK(clk), .RN(n469), .Q(
        fb_addr[5]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[4]  ( .D(n16), .CK(clk), .RN(n546), .Q(
        fb_addr[4]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[2]  ( .D(n18), .CK(clk), .RN(n469), .Q(
        fb_addr[2]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[0]  ( .D(n416), .CK(clk), .RN(n546), .Q(
        fb_addr[0]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[1]  ( .D(n20), .CK(clk), .RN(n546), .Q(
        fb_addr[1]) );
  DFFRX1 \data_path/si_reg/q_reg[11]  ( .D(n396), .CK(clk), .RN(n546), .Q(
        \data_path/si_w[11] ), .QN(n712) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[14]  ( .D(n386), .CK(clk), .RN(n469), 
        .Q(fb_addr[14]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[9]  ( .D(n401), .CK(clk), .RN(n546), .Q(
        fb_addr[9]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[10]  ( .D(n398), .CK(clk), .RN(n546), 
        .Q(fb_addr[10]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[8]  ( .D(n14), .CK(clk), .RN(n546), .Q(
        fb_addr[8]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[7]  ( .D(n404), .CK(clk), .RN(n546), .Q(
        fb_addr[7]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[3]  ( .D(n413), .CK(clk), .RN(n469), .Q(
        fb_addr[3]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[13]  ( .D(n389), .CK(clk), .RN(n469), 
        .Q(fb_addr[13]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[11]  ( .D(n395), .CK(clk), .RN(n546), 
        .Q(fb_addr[11]) );
  DFFRX1 \data_path/init_time_reg/q_reg[5]  ( .D(n334), .CK(clk), .RN(n469), 
        .Q(curr_time[5]) );
  DFFRX1 \data_path/init_time_reg/q_reg[8]  ( .D(n331), .CK(clk), .RN(n546), 
        .Q(curr_time[8]) );
  DFFRX1 \data_path/so_reg/q_reg[1]  ( .D(n365), .CK(clk), .RN(n469), .QN(n479) );
  DFFRX1 \data_path/so_reg/q_reg[22]  ( .D(n344), .CK(clk), .RN(n469), .Q(n781) );
  DFFRX1 \data_path/so_reg/q_reg[21]  ( .D(n345), .CK(clk), .RN(n469), .QN(
        n477) );
  DFFRX1 \data_path/so_reg/q_reg[15]  ( .D(n351), .CK(clk), .RN(n469), .QN(
        n486) );
  DFFRX1 \data_path/so_reg/q_reg[14]  ( .D(n352), .CK(clk), .RN(n469), .QN(
        n488) );
  DFFRX1 \data_path/so_reg/q_reg[5]  ( .D(n361), .CK(clk), .RN(n469), .QN(n492) );
  DFFRX1 \data_path/so_reg/q_reg[4]  ( .D(n362), .CK(clk), .RN(n469), .QN(n490) );
  DFFRX1 \data_path/so_reg/q_reg[3]  ( .D(n363), .CK(clk), .RN(n469), .QN(n484) );
  DFFRX1 \data_path/so_reg/q_reg[2]  ( .D(n364), .CK(clk), .RN(n469), .QN(n482) );
  DFFRX1 \data_path/so_reg/q_reg[29]  ( .D(n337), .CK(clk), .RN(n546), .Q(
        im_d_w[29]) );
  DFFRX1 \data_path/so_reg/q_reg[19]  ( .D(n347), .CK(clk), .RN(n469), .Q(
        im_d_w_19) );
  DFFRX1 \data_path/so_reg/q_reg[9]  ( .D(n357), .CK(clk), .RN(n469), .Q(
        im_d_w_9) );
  DFFRX1 \data_path/so_reg/q_reg[16]  ( .D(n350), .CK(clk), .RN(n469), .QN(
        n475) );
  DFFRX1 \data_path/so_reg/q_reg[6]  ( .D(n360), .CK(clk), .RN(n469), .QN(n494) );
  DFFRX1 \data_path/so_reg/q_reg[17]  ( .D(n349), .CK(clk), .RN(n469), .QN(
        n496) );
  DFFRX1 \data_path/so_reg/q_reg[7]  ( .D(n359), .CK(clk), .RN(n469), .QN(n498) );
  BUFX4 U435 ( .A(n731), .Y(n544) );
  CLKBUFX3 U436 ( .A(n732), .Y(n545) );
  AOI22XL U437 ( .A0(\intadd_1/SUM[0] ), .A1(n542), .B0(\intadd_1/SUM[1] ), 
        .B1(n541), .Y(n421) );
  OAI21XL U438 ( .A0(\data_path/si_w[8] ), .A1(n620), .B0(en_so), .Y(n422) );
  OAI21XL U439 ( .A0(n786), .A1(n729), .B0(n465), .Y(n423) );
  AOI22X1 U440 ( .A0(n786), .A1(n422), .B0(\data_path/si_w[8] ), .B1(n423), 
        .Y(n424) );
  NAND3X1 U441 ( .A(n421), .B(n646), .C(n424), .Y(n356) );
  AOI22XL U442 ( .A0(\intadd_2/SUM[0] ), .A1(n542), .B0(\intadd_2/SUM[1] ), 
        .B1(n541), .Y(n425) );
  OAI21XL U443 ( .A0(\data_path/si_w[0] ), .A1(n620), .B0(en_so), .Y(n426) );
  OAI21XL U444 ( .A0(n787), .A1(n729), .B0(n465), .Y(n427) );
  AOI22X1 U445 ( .A0(n787), .A1(n426), .B0(\data_path/si_w[0] ), .B1(n427), 
        .Y(n428) );
  NAND3X1 U446 ( .A(n425), .B(n646), .C(n428), .Y(n366) );
  AOI22XL U447 ( .A0(\intadd_0/SUM[0] ), .A1(n542), .B0(\intadd_0/SUM[1] ), 
        .B1(n541), .Y(n429) );
  OAI21XL U448 ( .A0(\data_path/si_w[16] ), .A1(n620), .B0(en_so), .Y(n430) );
  OAI21XL U449 ( .A0(n782), .A1(n729), .B0(n465), .Y(n431) );
  AOI22X1 U450 ( .A0(n782), .A1(n430), .B0(\data_path/si_w[16] ), .B1(n431), 
        .Y(n432) );
  NAND3X1 U451 ( .A(n429), .B(n646), .C(n432), .Y(n346) );
  NOR2X1 U452 ( .A(n643), .B(n694), .Y(n433) );
  OAI2BB2XL U453 ( .B0(n465), .B1(n514), .A0N(\intadd_0/SUM[6] ), .A1N(n543), 
        .Y(n434) );
  AOI211X1 U454 ( .A0(n776), .A1(n728), .B0(n433), .C0(n434), .Y(n435) );
  OAI211X1 U455 ( .A0(n727), .A1(n693), .B0(n646), .C0(n435), .Y(n339) );
  NOR4X1 U456 ( .A(\data_path/si_w[16] ), .B(\data_path/si_w[17] ), .C(
        \data_path/si_w[18] ), .D(\data_path/si_w[19] ), .Y(n436) );
  NOR4X1 U457 ( .A(\data_path/si_w[1] ), .B(\data_path/si_w[2] ), .C(
        \data_path/si_w[15] ), .D(\data_path/si_w[23] ), .Y(n437) );
  NOR4X1 U458 ( .A(\data_path/si_w[20] ), .B(\data_path/si_w[14] ), .C(
        \data_path/si_w[21] ), .D(\data_path/si_w[22] ), .Y(n438) );
  AND4X1 U459 ( .A(n437), .B(n438), .C(n522), .D(en_curr_photo_size), .Y(n439)
         );
  AND4X1 U460 ( .A(n501), .B(n436), .C(n508), .D(n439), .Y(n552) );
  AO22X1 U461 ( .A0(n541), .A1(\intadd_1/SUM[2] ), .B0(\intadd_1/SUM[1] ), 
        .B1(n542), .Y(n440) );
  AOI211X1 U462 ( .A0(n728), .A1(n785), .B0(n638), .C0(n440), .Y(n441) );
  NAND2X1 U463 ( .A(\intadd_1/SUM[0] ), .B(n543), .Y(n442) );
  OAI211X1 U464 ( .A0(n465), .A1(n523), .B0(n441), .C0(n442), .Y(n355) );
  CLKBUFX8 U465 ( .A(n546), .Y(n469) );
  AOI211X1 U466 ( .A0(curr_time[13]), .A1(n670), .B0(curr_time[15]), .C0(
        curr_time[14]), .Y(n677) );
  CLKBUFX8 U467 ( .A(n22), .Y(n546) );
  INVX16 U468 ( .A(n443), .Y(IM_D[9]) );
  INVX16 U469 ( .A(n445), .Y(IM_D[10]) );
  INVX16 U470 ( .A(n447), .Y(IM_D[11]) );
  INVX16 U471 ( .A(n449), .Y(IM_D[19]) );
  INVX16 U472 ( .A(n451), .Y(IM_D[20]) );
  INVX16 U473 ( .A(n453), .Y(IM_D[21]) );
  INVX16 U474 ( .A(n455), .Y(IM_D[22]) );
  INVX16 U475 ( .A(n457), .Y(IM_D[23]) );
  INVX16 U476 ( .A(n459), .Y(IM_D[8]) );
  INVX16 U477 ( .A(n461), .Y(IM_D[0]) );
  INVX16 U478 ( .A(n463), .Y(IM_D[16]) );
  INVX12 U479 ( .A(reset), .Y(n22) );
  BUFX4 U480 ( .A(n645), .Y(n465) );
  NOR2X1 U481 ( .A(n658), .B(n660), .Y(n666) );
  INVX6 U482 ( .A(n548), .Y(n466) );
  INVX6 U483 ( .A(n547), .Y(n467) );
  INVX6 U484 ( .A(en_so), .Y(n728) );
  INVX3 U485 ( .A(en_si), .Y(n732) );
  NOR2X2 U486 ( .A(expand_sel[1]), .B(expand_sel[0]), .Y(n571) );
  CLKINVX1 U487 ( .A(n468), .Y(n547) );
  NOR2X1 U488 ( .A(si_sel), .B(n545), .Y(n731) );
  INVX16 U489 ( .A(n486), .Y(IM_D[13]) );
  BUFX16 U490 ( .A(n781), .Y(IM_D[18]) );
  NAND2X1 U491 ( .A(n710), .B(n709), .Y(n720) );
  NOR2X1 U492 ( .A(n506), .B(n708), .Y(n709) );
  NOR2X1 U493 ( .A(n531), .B(n658), .Y(n661) );
  NAND2X1 U494 ( .A(curr_time[2]), .B(n655), .Y(n658) );
  NOR2X1 U495 ( .A(n699), .B(n724), .Y(n703) );
  NOR2X1 U496 ( .A(curr_time[8]), .B(n715), .Y(n699) );
  CLKINVX1 U497 ( .A(n649), .Y(n660) );
  NOR2X1 U498 ( .A(n671), .B(n664), .Y(n649) );
  NOR2X1 U499 ( .A(n503), .B(n686), .Y(n681) );
  NAND2X1 U500 ( .A(en_init_time), .B(n679), .Y(n686) );
  AOI211X1 U501 ( .A0(n647), .A1(curr_time[5]), .B0(curr_time[6]), .C0(
        curr_time[7]), .Y(n669) );
  OAI21X1 U502 ( .A0(curr_time[16]), .A1(n687), .B0(n722), .Y(n682) );
  CLKINVX1 U503 ( .A(n679), .Y(n687) );
  AOI211X1 U504 ( .A0(n688), .A1(curr_time[20]), .B0(n677), .C0(n676), .Y(n679) );
  NOR2BX1 U505 ( .AN(init_time_mux_sel), .B(n669), .Y(n675) );
  AOI211X1 U506 ( .A0(curr_time[2]), .A1(n655), .B0(n671), .C0(n664), .Y(n656)
         );
  NAND2X1 U507 ( .A(n669), .B(init_time_mux_sel), .Y(n664) );
  NOR2BX1 U508 ( .AN(n688), .B(n686), .Y(n690) );
  OAI21X1 U509 ( .A0(n688), .A1(n687), .B0(n722), .Y(n691) );
  NOR3X2 U510 ( .A(n507), .B(n503), .C(n521), .Y(n688) );
  OAI21X1 U511 ( .A0(\intadd_0/n1 ), .A1(im_d_w[28]), .B0(n642), .Y(n693) );
  NAND2X1 U512 ( .A(\intadd_0/n1 ), .B(im_d_w[28]), .Y(n642) );
  OAI31X1 U513 ( .A0(n562), .A1(n561), .A2(n560), .B0(expand_sel[3]), .Y(n576)
         );
  CLKINVX1 U514 ( .A(n541), .Y(n643) );
  BUFX4 U515 ( .A(n633), .Y(n541) );
  BUFX4 U516 ( .A(n639), .Y(n542) );
  CLKINVX1 U517 ( .A(n736), .Y(n471) );
  INVX16 U518 ( .A(n471), .Y(IM_A[0]) );
  INVX16 U519 ( .A(n774), .Y(IM_A[1]) );
  INVX16 U520 ( .A(n773), .Y(IM_A[2]) );
  INVX16 U521 ( .A(n772), .Y(IM_A[3]) );
  INVX16 U522 ( .A(n771), .Y(IM_A[4]) );
  INVX16 U523 ( .A(n770), .Y(IM_A[5]) );
  INVX16 U524 ( .A(n769), .Y(IM_A[6]) );
  INVX16 U525 ( .A(n768), .Y(IM_A[7]) );
  INVX16 U526 ( .A(n767), .Y(IM_A[8]) );
  INVX16 U527 ( .A(n766), .Y(IM_A[9]) );
  INVX16 U528 ( .A(n765), .Y(IM_A[10]) );
  INVX16 U529 ( .A(n764), .Y(IM_A[11]) );
  INVX16 U530 ( .A(n763), .Y(IM_A[12]) );
  INVX16 U531 ( .A(n762), .Y(IM_A[13]) );
  INVX16 U532 ( .A(n761), .Y(IM_A[14]) );
  INVX16 U533 ( .A(n760), .Y(IM_A[15]) );
  INVX16 U534 ( .A(n759), .Y(IM_A[16]) );
  INVX16 U535 ( .A(n758), .Y(IM_A[17]) );
  INVX16 U536 ( .A(n757), .Y(IM_A[18]) );
  CLKINVX1 U537 ( .A(n755), .Y(n473) );
  INVX16 U538 ( .A(n473), .Y(IM_A[19]) );
  INVX16 U539 ( .A(n475), .Y(IM_D[14]) );
  INVX16 U540 ( .A(n477), .Y(IM_D[17]) );
  INVX16 U541 ( .A(n479), .Y(IM_D[1]) );
  INVX16 U542 ( .A(n482), .Y(IM_D[2]) );
  INVX16 U543 ( .A(n484), .Y(IM_D[3]) );
  INVX16 U544 ( .A(n488), .Y(IM_D[12]) );
  INVX16 U545 ( .A(n490), .Y(IM_D[4]) );
  INVX16 U546 ( .A(n492), .Y(IM_D[5]) );
  INVX16 U547 ( .A(n494), .Y(IM_D[6]) );
  INVX16 U548 ( .A(n496), .Y(IM_D[15]) );
  INVX16 U549 ( .A(n498), .Y(IM_D[7]) );
  NAND2X1 U550 ( .A(expand_sel[0]), .B(n568), .Y(n569) );
  NOR2X1 U551 ( .A(curr_time[2]), .B(n655), .Y(n653) );
  NOR2X2 U552 ( .A(n650), .B(n517), .Y(n655) );
  OAI21X1 U553 ( .A0(\intadd_2/n1 ), .A1(im_d_w_8), .B0(n596), .Y(n600) );
  NAND2X1 U554 ( .A(\intadd_2/n1 ), .B(im_d_w_8), .Y(n596) );
  OAI21X1 U555 ( .A0(\intadd_1/n1 ), .A1(im_d_w_18), .B0(n616), .Y(n726) );
  NAND2X1 U556 ( .A(\intadd_1/n1 ), .B(im_d_w_18), .Y(n616) );
  NOR2X1 U557 ( .A(\data_path/si_w[4] ), .B(n550), .Y(n553) );
  NAND4X1 U558 ( .A(n500), .B(n712), .C(n509), .D(n524), .Y(n550) );
  NAND2X1 U559 ( .A(n557), .B(n470), .Y(n620) );
  CLKINVX1 U560 ( .A(n710), .Y(n715) );
  NOR2X1 U561 ( .A(n673), .B(n671), .Y(n710) );
  CLKINVX1 U562 ( .A(expand_sel[1]), .Y(n568) );
  NAND2XL U563 ( .A(IM_D[14]), .B(n728), .Y(n614) );
  BUFX4 U564 ( .A(n644), .Y(n543) );
  NOR2XL U565 ( .A(n728), .B(n620), .Y(n644) );
  INVX3 U566 ( .A(n725), .Y(n723) );
  NOR2X4 U567 ( .A(init_time_mux_sel), .B(n671), .Y(n725) );
  INVX4 U568 ( .A(n646), .Y(n638) );
  NAND4X2 U569 ( .A(\so_mux_sel[1] ), .B(n577), .C(n576), .D(n575), .Y(n646)
         );
  NOR2BX2 U570 ( .AN(n673), .B(n724), .Y(n722) );
  NAND2X2 U571 ( .A(en_init_time), .B(n664), .Y(n724) );
  NAND2XL U572 ( .A(n777), .B(n728), .Y(n640) );
  INVXL U573 ( .A(en_photo_num), .Y(n734) );
  OAI211XL U574 ( .A0(en_curr_photo_size), .A1(n515), .B0(n555), .C0(n735), 
        .Y(n368) );
  NAND4XL U575 ( .A(\data_path/si_w[7] ), .B(n553), .C(n552), .D(n551), .Y(
        n555) );
  NOR3XL U576 ( .A(\data_path/si_w[9] ), .B(\data_path/si_w[0] ), .C(
        \data_path/si_w[3] ), .Y(n551) );
  NAND4XL U577 ( .A(n554), .B(n553), .C(n552), .D(n519), .Y(n735) );
  INVXL U578 ( .A(n702), .Y(n402) );
  INVXL U579 ( .A(n696), .Y(n411) );
  INVXL U580 ( .A(n707), .Y(n399) );
  INVXL U581 ( .A(n695), .Y(n414) );
  INVXL U582 ( .A(n698), .Y(n405) );
  INVXL U583 ( .A(n719), .Y(n393) );
  INVXL U584 ( .A(n713), .Y(n396) );
  INVXL U585 ( .A(n697), .Y(n408) );
  INVXL U586 ( .A(n653), .Y(n654) );
  AOI211XL U587 ( .A0(curr_time[4]), .A1(n671), .B0(n663), .C0(n662), .Y(n141)
         );
  NOR2XL U588 ( .A(n723), .B(n510), .Y(n662) );
  AOI211XL U589 ( .A0(curr_time[4]), .A1(n661), .B0(n660), .C0(n659), .Y(n663)
         );
  NOR2XL U590 ( .A(curr_time[4]), .B(n661), .Y(n659) );
  NOR2XL U591 ( .A(n652), .B(n651), .Y(n145) );
  AOI211XL U592 ( .A0(n650), .A1(n517), .B0(n655), .C0(n660), .Y(n652) );
  INVXL U593 ( .A(n668), .Y(n334) );
  INVXL U594 ( .A(n665), .Y(n667) );
  OAI32XL U595 ( .A0(n531), .A1(n656), .A2(n671), .B0(n666), .B1(curr_time[3]), 
        .Y(n657) );
  AOI21XL U596 ( .A0(curr_time[8]), .A1(n724), .B0(n699), .Y(n672) );
  NAND2XL U597 ( .A(curr_time[12]), .B(curr_time[11]), .Y(n721) );
  AOI22XL U598 ( .A0(curr_time[12]), .A1(n716), .B0(n725), .B1(
        \data_path/si_w[12] ), .Y(n717) );
  AOI22XL U599 ( .A0(curr_time[10]), .A1(n704), .B0(\data_path/si_w[10] ), 
        .B1(n725), .Y(n705) );
  NAND2XL U600 ( .A(curr_time[8]), .B(n710), .Y(n706) );
  OAI211XL U601 ( .A0(n723), .A1(n526), .B0(n685), .C0(n684), .Y(n321) );
  NOR2XL U602 ( .A(n687), .B(curr_time[17]), .Y(n683) );
  NAND3XL U603 ( .A(curr_time[17]), .B(n681), .C(n521), .Y(n685) );
  INVXL U604 ( .A(n692), .Y(n319) );
  NAND2XL U605 ( .A(n675), .B(n677), .Y(n673) );
  NAND3XL U606 ( .A(n675), .B(n674), .C(n504), .Y(n676) );
  AOI211XL U607 ( .A0(curr_time[20]), .A1(curr_time[19]), .B0(curr_time[21]), 
        .C0(curr_time[22]), .Y(n674) );
  NOR2XL U608 ( .A(n653), .B(n665), .Y(n647) );
  NAND2XL U609 ( .A(curr_time[4]), .B(curr_time[3]), .Y(n665) );
  AOI211XL U610 ( .A0(n506), .A1(n708), .B0(n520), .C0(n502), .Y(n670) );
  NAND2XL U611 ( .A(curr_time[9]), .B(curr_time[8]), .Y(n708) );
  CLKINVX2 U612 ( .A(en_init_time), .Y(n671) );
  OAI211XL U613 ( .A0(n465), .A1(n509), .B0(n592), .C0(n591), .Y(n361) );
  NAND2XL U614 ( .A(n543), .B(\intadd_2/SUM[4] ), .Y(n591) );
  AOI211XL U615 ( .A0(n542), .A1(\intadd_2/SUM[5] ), .B0(n638), .C0(n590), .Y(
        n592) );
  OAI211XL U616 ( .A0(n512), .A1(n465), .B0(n636), .C0(n635), .Y(n341) );
  NAND2XL U617 ( .A(n543), .B(\intadd_0/SUM[4] ), .Y(n635) );
  AOI211XL U618 ( .A0(n542), .A1(\intadd_0/SUM[5] ), .B0(n638), .C0(n634), .Y(
        n636) );
  OAI211XL U619 ( .A0(n465), .A1(n527), .B0(n623), .C0(n622), .Y(n345) );
  NAND2XL U620 ( .A(n543), .B(\intadd_0/SUM[0] ), .Y(n622) );
  AOI211XL U621 ( .A0(n542), .A1(\intadd_0/SUM[1] ), .B0(n638), .C0(n621), .Y(
        n623) );
  OAI211XL U622 ( .A0(n465), .A1(n522), .B0(n609), .C0(n608), .Y(n352) );
  NAND2XL U623 ( .A(n543), .B(\intadd_1/SUM[3] ), .Y(n608) );
  AOI211XL U624 ( .A0(n542), .A1(\intadd_1/SUM[4] ), .B0(n638), .C0(n607), .Y(
        n609) );
  OAI211XL U625 ( .A0(n465), .A1(n510), .B0(n589), .C0(n588), .Y(n362) );
  NAND2XL U626 ( .A(n543), .B(\intadd_2/SUM[3] ), .Y(n588) );
  AOI211XL U627 ( .A0(n542), .A1(\intadd_2/SUM[4] ), .B0(n638), .C0(n587), .Y(
        n589) );
  OAI211XL U628 ( .A0(n465), .A1(n500), .B0(n603), .C0(n602), .Y(n354) );
  NAND2XL U629 ( .A(n543), .B(\intadd_1/SUM[1] ), .Y(n602) );
  AOI211XL U630 ( .A0(n542), .A1(\intadd_1/SUM[2] ), .B0(n638), .C0(n601), .Y(
        n603) );
  OAI211XL U631 ( .A0(n465), .A1(n712), .B0(n606), .C0(n605), .Y(n353) );
  NAND2XL U632 ( .A(n543), .B(\intadd_1/SUM[2] ), .Y(n605) );
  AOI211XL U633 ( .A0(n542), .A1(\intadd_1/SUM[3] ), .B0(n638), .C0(n604), .Y(
        n606) );
  OAI211XL U634 ( .A0(n465), .A1(n528), .B0(n629), .C0(n628), .Y(n343) );
  NAND2XL U635 ( .A(n543), .B(\intadd_0/SUM[2] ), .Y(n628) );
  AOI211XL U636 ( .A0(n542), .A1(\intadd_0/SUM[3] ), .B0(n638), .C0(n627), .Y(
        n629) );
  OAI211XL U637 ( .A0(n465), .A1(n518), .B0(n586), .C0(n585), .Y(n363) );
  NAND2XL U638 ( .A(n543), .B(\intadd_2/SUM[2] ), .Y(n585) );
  AOI211XL U639 ( .A0(n542), .A1(\intadd_2/SUM[3] ), .B0(n638), .C0(n584), .Y(
        n586) );
  OAI211XL U640 ( .A0(n508), .A1(n465), .B0(n612), .C0(n611), .Y(n351) );
  NAND2XL U641 ( .A(n543), .B(\intadd_1/SUM[4] ), .Y(n611) );
  AOI211XL U642 ( .A0(n542), .A1(\intadd_1/SUM[5] ), .B0(n638), .C0(n610), .Y(
        n612) );
  OAI211XL U643 ( .A0(n465), .A1(n505), .B0(n580), .C0(n579), .Y(n365) );
  NAND2XL U644 ( .A(n543), .B(\intadd_2/SUM[0] ), .Y(n579) );
  AOI211XL U645 ( .A0(\intadd_2/SUM[1] ), .A1(n542), .B0(n638), .C0(n578), .Y(
        n580) );
  OAI211XL U646 ( .A0(n465), .A1(n511), .B0(n583), .C0(n582), .Y(n364) );
  NAND2XL U647 ( .A(n543), .B(\intadd_2/SUM[1] ), .Y(n582) );
  AOI211XL U648 ( .A0(n542), .A1(\intadd_2/SUM[2] ), .B0(n638), .C0(n581), .Y(
        n583) );
  OAI211XL U649 ( .A0(n465), .A1(n534), .B0(n632), .C0(n631), .Y(n342) );
  NAND2XL U650 ( .A(n543), .B(\intadd_0/SUM[3] ), .Y(n631) );
  AOI211XL U651 ( .A0(n542), .A1(\intadd_0/SUM[4] ), .B0(n638), .C0(n630), .Y(
        n632) );
  OAI211XL U652 ( .A0(n465), .A1(n526), .B0(n626), .C0(n625), .Y(n344) );
  NAND2XL U653 ( .A(n543), .B(\intadd_0/SUM[1] ), .Y(n625) );
  AOI211XL U654 ( .A0(n542), .A1(\intadd_0/SUM[2] ), .B0(n638), .C0(n624), .Y(
        n626) );
  OAI211XL U655 ( .A0(n693), .A1(n643), .B0(n641), .C0(n640), .Y(n340) );
  AOI211XL U656 ( .A0(n542), .A1(\intadd_0/SUM[6] ), .B0(n638), .C0(n637), .Y(
        n641) );
  OAI211XL U657 ( .A0(n600), .A1(n643), .B0(n595), .C0(n594), .Y(n360) );
  NAND2X1 U658 ( .A(IM_D[6]), .B(n728), .Y(n594) );
  AOI211XL U659 ( .A0(n542), .A1(\intadd_2/SUM[6] ), .B0(n638), .C0(n593), .Y(
        n595) );
  OAI211XL U660 ( .A0(n726), .A1(n643), .B0(n615), .C0(n614), .Y(n350) );
  AOI211XL U661 ( .A0(n542), .A1(\intadd_1/SUM[6] ), .B0(n638), .C0(n613), .Y(
        n615) );
  OAI211XL U662 ( .A0(n727), .A1(n600), .B0(n599), .C0(n646), .Y(n359) );
  AOI211X1 U663 ( .A0(IM_D[7]), .A1(n728), .B0(n598), .C0(n597), .Y(n599) );
  NOR2XL U664 ( .A(n643), .B(n701), .Y(n598) );
  OAI211XL U665 ( .A0(n727), .A1(n726), .B0(n619), .C0(n646), .Y(n349) );
  AOI211X1 U666 ( .A0(IM_D[15]), .A1(n728), .B0(n618), .C0(n617), .Y(n619) );
  NOR2XL U667 ( .A(n643), .B(n730), .Y(n618) );
  AND2XL U668 ( .A(\data_path/si_w[16] ), .B(n782), .Y(\intadd_0/CI ) );
  NOR2BXL U669 ( .AN(n787), .B(n516), .Y(\intadd_2/CI ) );
  INVXL U670 ( .A(expand_sel[3]), .Y(n572) );
  AOI211XL U671 ( .A0(n571), .A1(\data_path/si_w[12] ), .B0(expand_sel[2]), 
        .C0(n570), .Y(n573) );
  AOI211XL U672 ( .A0(n571), .A1(\data_path/si_w[8] ), .B0(n565), .C0(n564), 
        .Y(n574) );
  AOI211XL U673 ( .A0(n571), .A1(\data_path/si_w[4] ), .B0(expand_sel[2]), 
        .C0(n559), .Y(n560) );
  INVXL U674 ( .A(expand_sel[0]), .Y(n566) );
  NOR2XL U675 ( .A(\data_path/si_w[0] ), .B(n565), .Y(n561) );
  NOR2XL U676 ( .A(n571), .B(n565), .Y(n562) );
  INVXL U677 ( .A(expand_sel[2]), .Y(n565) );
  NOR2XL U678 ( .A(n470), .B(n728), .Y(n577) );
  INVX3 U679 ( .A(n543), .Y(n729) );
  INVXL U680 ( .A(\so_mux_sel[1] ), .Y(n557) );
  NOR2BXL U681 ( .AN(n786), .B(n501), .Y(\intadd_1/CI ) );
  NOR2BXL U682 ( .AN(\sftr_n[1] ), .B(n556), .Y(n633) );
  NAND3XL U683 ( .A(\so_mux_sel[1] ), .B(n470), .C(en_so), .Y(n556) );
  INVXL U684 ( .A(n775), .Y(n736) );
  INVXL U685 ( .A(n756), .Y(n755) );
  OAI22XL U686 ( .A0(en_photo_num), .A1(n10), .B0(n734), .B1(n733), .Y(n21) );
  AOI222XL U687 ( .A0(n732), .A1(\data_path/si_w[2] ), .B0(n544), .B1(IM_Q[2]), 
        .C0(n718), .C1(CR_Q[2]), .Y(n314) );
  AOI222XL U688 ( .A0(n545), .A1(\data_path/si_w[8] ), .B0(n544), .B1(IM_Q[8]), 
        .C0(n718), .C1(CR_Q[8]), .Y(n312) );
  AOI222XL U689 ( .A0(n545), .A1(\data_path/si_w[4] ), .B0(n544), .B1(IM_Q[4]), 
        .C0(n718), .C1(CR_Q[4]), .Y(n313) );
  AOI222XL U690 ( .A0(n545), .A1(\data_path/si_w[1] ), .B0(n718), .B1(CR_Q[1]), 
        .C0(IM_Q[1]), .C1(n544), .Y(n315) );
  NOR3XL U691 ( .A(\data_path/si_w[0] ), .B(\data_path/si_w[3] ), .C(n523), 
        .Y(n554) );
  AOI222XL U692 ( .A0(n545), .A1(\data_path/si_w[9] ), .B0(n544), .B1(IM_Q[9]), 
        .C0(n718), .C1(CR_Q[9]), .Y(n702) );
  AOI222XL U693 ( .A0(n545), .A1(\data_path/si_w[5] ), .B0(n544), .B1(IM_Q[5]), 
        .C0(n718), .C1(CR_Q[5]), .Y(n696) );
  AOI222XL U694 ( .A0(n545), .A1(\data_path/si_w[0] ), .B0(n544), .B1(IM_Q[0]), 
        .C0(n718), .C1(CR_Q[0]), .Y(n549) );
  CLKINVX1 U695 ( .A(en_fb_addr), .Y(n548) );
  AOI222XL U696 ( .A0(n545), .A1(\data_path/si_w[10] ), .B0(n544), .B1(
        IM_Q[10]), .C0(n718), .C1(CR_Q[10]), .Y(n707) );
  AOI222XL U697 ( .A0(n545), .A1(\data_path/si_w[3] ), .B0(n544), .B1(IM_Q[3]), 
        .C0(n718), .C1(CR_Q[3]), .Y(n695) );
  AOI222XL U698 ( .A0(n545), .A1(\data_path/si_w[7] ), .B0(n544), .B1(IM_Q[7]), 
        .C0(n718), .C1(CR_Q[7]), .Y(n698) );
  AOI222XL U699 ( .A0(n545), .A1(\data_path/si_w[12] ), .B0(n544), .B1(
        IM_Q[12]), .C0(n718), .C1(CR_Q[12]), .Y(n719) );
  AOI222XL U700 ( .A0(n545), .A1(\data_path/si_w[11] ), .B0(n544), .B1(
        IM_Q[11]), .C0(n718), .C1(CR_Q[11]), .Y(n713) );
  AOI222XL U701 ( .A0(n545), .A1(\data_path/si_w[6] ), .B0(n544), .B1(IM_Q[6]), 
        .C0(n718), .C1(CR_Q[6]), .Y(n697) );
  AND2X2 U702 ( .A(si_sel), .B(en_si), .Y(n718) );
  AOI222XL U703 ( .A0(n671), .A1(curr_time[2]), .B0(n725), .B1(
        \data_path/si_w[2] ), .C0(n654), .C1(n656), .Y(n144) );
  AOI222XL U704 ( .A0(\data_path/si_w[5] ), .A1(n725), .B0(curr_time[5]), .B1(
        n724), .C0(n667), .C1(n666), .Y(n668) );
  OAI21XL U705 ( .A0(n714), .A1(n502), .B0(n711), .Y(n328) );
  OAI222XL U706 ( .A0(n508), .A1(n723), .B0(n535), .B1(n722), .C0(n721), .C1(
        n720), .Y(n326) );
  OAI31XL U707 ( .A0(curr_time[12]), .A1(n502), .A2(n720), .B0(n717), .Y(n327)
         );
  OAI31XL U708 ( .A0(curr_time[10]), .A1(n530), .A2(n706), .B0(n705), .Y(n329)
         );
  AOI222XL U709 ( .A0(n691), .A1(curr_time[20]), .B0(curr_time[19]), .B1(n690), 
        .C0(n725), .C1(\data_path/si_w[20] ), .Y(n692) );
  CLKINVX1 U710 ( .A(n542), .Y(n727) );
  NAND3BX1 U711 ( .AN(n470), .B(en_so), .C(n557), .Y(n645) );
  NOR2X1 U712 ( .A(\sftr_n[1] ), .B(n556), .Y(n639) );
  AO22X1 U713 ( .A0(\data_path/si_w[16] ), .A1(n732), .B0(n544), .B1(IM_Q[16]), 
        .Y(n418) );
  AOI2BB2X1 U714 ( .B0(n466), .B1(n516), .A0N(en_fb_addr), .A1N(fb_addr[0]), 
        .Y(n416) );
  AOI2BB2X1 U715 ( .B0(n467), .B1(n516), .A0N(n467), .A1N(curr_photo_addr[0]), 
        .Y(n415) );
  AOI2BB2X1 U716 ( .B0(n466), .B1(n518), .A0N(n466), .A1N(fb_addr[3]), .Y(n413) );
  AOI2BB2X1 U717 ( .B0(n467), .B1(n518), .A0N(n467), .A1N(curr_photo_addr[3]), 
        .Y(n412) );
  AOI2BB2X1 U718 ( .B0(n466), .B1(n509), .A0N(en_fb_addr), .A1N(fb_addr[5]), 
        .Y(n410) );
  AOI2BB2X1 U719 ( .B0(n467), .B1(n509), .A0N(n467), .A1N(curr_photo_addr[5]), 
        .Y(n409) );
  AOI2BB2X1 U720 ( .B0(n466), .B1(n524), .A0N(en_fb_addr), .A1N(fb_addr[6]), 
        .Y(n407) );
  AOI2BB2X1 U721 ( .B0(n467), .B1(n524), .A0N(n467), .A1N(curr_photo_addr[6]), 
        .Y(n406) );
  AOI2BB2X1 U722 ( .B0(n466), .B1(n519), .A0N(n466), .A1N(fb_addr[7]), .Y(n404) );
  AOI2BB2X1 U723 ( .B0(n467), .B1(n519), .A0N(n467), .A1N(curr_photo_addr[7]), 
        .Y(n403) );
  AOI2BB2X1 U724 ( .B0(en_photo_num), .B1(\data_path/si_w[0] ), .A0N(
        en_photo_num), .A1N(photo_num[0]), .Y(n367) );
  OAI22XL U725 ( .A0(expand_sel[0]), .A1(\data_path/si_w[2] ), .B0(n566), .B1(
        \data_path/si_w[1] ), .Y(n558) );
  OAI22XL U726 ( .A0(n568), .A1(n558), .B0(n518), .B1(n569), .Y(n559) );
  OAI22XL U727 ( .A0(expand_sel[0]), .A1(\data_path/si_w[6] ), .B0(n566), .B1(
        \data_path/si_w[5] ), .Y(n563) );
  OAI22XL U728 ( .A0(n568), .A1(n563), .B0(n569), .B1(n519), .Y(n564) );
  OAI22XL U729 ( .A0(expand_sel[0]), .A1(\data_path/si_w[10] ), .B0(n566), 
        .B1(\data_path/si_w[9] ), .Y(n567) );
  OAI22XL U730 ( .A0(n712), .A1(n569), .B0(n568), .B1(n567), .Y(n570) );
  OAI21XL U731 ( .A0(n574), .A1(n573), .B0(n572), .Y(n575) );
  AO22X1 U732 ( .A0(\intadd_2/SUM[2] ), .A1(n541), .B0(IM_D[1]), .B1(n728), 
        .Y(n578) );
  AO22X1 U733 ( .A0(\intadd_2/SUM[3] ), .A1(n541), .B0(IM_D[2]), .B1(n728), 
        .Y(n581) );
  AO22X1 U734 ( .A0(\intadd_2/SUM[4] ), .A1(n541), .B0(IM_D[3]), .B1(n728), 
        .Y(n584) );
  AO22X1 U735 ( .A0(\intadd_2/SUM[5] ), .A1(n541), .B0(IM_D[4]), .B1(n728), 
        .Y(n587) );
  AO22X1 U736 ( .A0(\intadd_2/SUM[6] ), .A1(n541), .B0(IM_D[5]), .B1(n728), 
        .Y(n590) );
  OAI2BB2XL U737 ( .B0(n524), .B1(n465), .A0N(n543), .A1N(\intadd_2/SUM[5] ), 
        .Y(n593) );
  AOI2BB2X1 U738 ( .B0(im_d_w_9), .B1(n596), .A0N(im_d_w_9), .A1N(n596), .Y(
        n701) );
  OAI2BB2XL U739 ( .B0(n519), .B1(n465), .A0N(n543), .A1N(\intadd_2/SUM[6] ), 
        .Y(n597) );
  OAI222XL U740 ( .A0(n701), .A1(n727), .B0(n538), .B1(en_so), .C0(n600), .C1(
        n729), .Y(n358) );
  AO22X1 U741 ( .A0(\intadd_1/SUM[3] ), .A1(n541), .B0(n784), .B1(n728), .Y(
        n601) );
  AO22X1 U742 ( .A0(\intadd_1/SUM[4] ), .A1(n541), .B0(n783), .B1(n728), .Y(
        n604) );
  AO22X1 U743 ( .A0(\intadd_1/SUM[5] ), .A1(n541), .B0(IM_D[12]), .B1(n728), 
        .Y(n607) );
  AO22X1 U744 ( .A0(\intadd_1/SUM[6] ), .A1(n541), .B0(IM_D[13]), .B1(n728), 
        .Y(n610) );
  OAI2BB2XL U745 ( .B0(n465), .B1(n529), .A0N(n543), .A1N(\intadd_1/SUM[5] ), 
        .Y(n613) );
  AOI2BB2X1 U746 ( .B0(im_d_w_19), .B1(n616), .A0N(im_d_w_19), .A1N(n616), .Y(
        n730) );
  OAI2BB2XL U747 ( .B0(n465), .B1(n525), .A0N(n543), .A1N(\intadd_1/SUM[6] ), 
        .Y(n617) );
  AO22X1 U748 ( .A0(\intadd_0/SUM[2] ), .A1(n541), .B0(IM_D[17]), .B1(n728), 
        .Y(n621) );
  AO22X1 U749 ( .A0(\intadd_0/SUM[3] ), .A1(n541), .B0(IM_D[18]), .B1(n728), 
        .Y(n624) );
  AO22X1 U750 ( .A0(\intadd_0/SUM[4] ), .A1(n541), .B0(n780), .B1(n728), .Y(
        n627) );
  AO22X1 U751 ( .A0(\intadd_0/SUM[5] ), .A1(n541), .B0(n779), .B1(n728), .Y(
        n630) );
  AO22X1 U752 ( .A0(\intadd_0/SUM[6] ), .A1(n541), .B0(n778), .B1(n728), .Y(
        n634) );
  OAI2BB2XL U753 ( .B0(n465), .B1(n513), .A0N(n543), .A1N(\intadd_0/SUM[5] ), 
        .Y(n637) );
  AOI2BB2X1 U754 ( .B0(im_d_w[29]), .B1(n642), .A0N(im_d_w[29]), .A1N(n642), 
        .Y(n694) );
  OAI22XL U755 ( .A0(curr_time[0]), .A1(n649), .B0(n517), .B1(n671), .Y(n648)
         );
  OAI21XL U756 ( .A0(n723), .A1(n516), .B0(n648), .Y(n336) );
  OAI22XL U757 ( .A0(en_init_time), .A1(n650), .B0(n723), .B1(n505), .Y(n651)
         );
  OAI21XL U758 ( .A0(n723), .A1(n518), .B0(n657), .Y(n335) );
  AO22X1 U759 ( .A0(n725), .A1(\data_path/si_w[6] ), .B0(n671), .B1(
        curr_time[6]), .Y(n333) );
  AO22X1 U760 ( .A0(n725), .A1(\data_path/si_w[7] ), .B0(n671), .B1(
        curr_time[7]), .Y(n332) );
  OAI21XL U761 ( .A0(n723), .A1(n501), .B0(n672), .Y(n331) );
  AOI2BB2X1 U762 ( .B0(n725), .B1(\data_path/si_w[16] ), .A0N(curr_time[16]), 
        .A1N(n686), .Y(n678) );
  OAI21XL U763 ( .A0(n722), .A1(n503), .B0(n678), .Y(n323) );
  OAI22XL U764 ( .A0(curr_time[17]), .A1(n681), .B0(n507), .B1(n682), .Y(n680)
         );
  OAI21XL U765 ( .A0(n723), .A1(n527), .B0(n680), .Y(n322) );
  OAI21XL U766 ( .A0(n683), .A1(n682), .B0(curr_time[18]), .Y(n684) );
  OAI22XL U767 ( .A0(curr_time[19]), .A1(n690), .B0(n533), .B1(n691), .Y(n689)
         );
  OAI21XL U768 ( .A0(n723), .A1(n528), .B0(n689), .Y(n320) );
  OAI22XL U769 ( .A0(n722), .A1(n536), .B0(n723), .B1(n512), .Y(n318) );
  OAI22XL U770 ( .A0(n722), .A1(n532), .B0(n723), .B1(n513), .Y(n317) );
  OAI22XL U771 ( .A0(n722), .A1(n504), .B0(n723), .B1(n514), .Y(n316) );
  OAI222XL U772 ( .A0(n694), .A1(n727), .B0(n539), .B1(en_so), .C0(n693), .C1(
        n729), .Y(n338) );
  OAI2BB2XL U773 ( .B0(n694), .B1(n729), .A0N(im_d_w[29]), .A1N(n728), .Y(n337) );
  AOI2BB2X1 U774 ( .B0(\data_path/si_w[9] ), .B1(n725), .A0N(curr_time[9]), 
        .A1N(n706), .Y(n700) );
  OAI21XL U775 ( .A0(n703), .A1(n530), .B0(n700), .Y(n330) );
  OAI2BB2XL U776 ( .B0(n701), .B1(n729), .A0N(im_d_w_9), .A1N(n728), .Y(n357)
         );
  AOI2BB2X1 U777 ( .B0(n467), .B1(n523), .A0N(n467), .A1N(curr_photo_addr[9]), 
        .Y(n400) );
  AOI2BB2X1 U778 ( .B0(n466), .B1(n523), .A0N(n466), .A1N(fb_addr[9]), .Y(n401) );
  OAI21XL U779 ( .A0(curr_time[9]), .A1(n715), .B0(n703), .Y(n704) );
  AOI2BB2X1 U780 ( .B0(n467), .B1(n500), .A0N(n467), .A1N(curr_photo_addr[10]), 
        .Y(n397) );
  AOI2BB2X1 U781 ( .B0(n466), .B1(n500), .A0N(n466), .A1N(fb_addr[10]), .Y(
        n398) );
  AOI2BB1X1 U782 ( .A0N(n709), .A1N(n715), .B0(n724), .Y(n714) );
  AOI2BB2X1 U783 ( .B0(\data_path/si_w[11] ), .B1(n725), .A0N(curr_time[11]), 
        .A1N(n720), .Y(n711) );
  AOI2BB2X1 U784 ( .B0(n467), .B1(n712), .A0N(n467), .A1N(curr_photo_addr[11]), 
        .Y(n394) );
  AOI2BB2X1 U785 ( .B0(n466), .B1(n712), .A0N(n466), .A1N(fb_addr[11]), .Y(
        n395) );
  OAI21XL U786 ( .A0(curr_time[11]), .A1(n715), .B0(n714), .Y(n716) );
  AOI2BB2X1 U787 ( .B0(n467), .B1(n522), .A0N(n467), .A1N(curr_photo_addr[12]), 
        .Y(n391) );
  AOI2BB2X1 U788 ( .B0(n466), .B1(n522), .A0N(en_fb_addr), .A1N(fb_addr[12]), 
        .Y(n392) );
  AOI2BB2X1 U789 ( .B0(n467), .B1(n508), .A0N(n467), .A1N(curr_photo_addr[13]), 
        .Y(n388) );
  AOI2BB2X1 U790 ( .B0(n466), .B1(n508), .A0N(n466), .A1N(fb_addr[13]), .Y(
        n389) );
  AO22X1 U791 ( .A0(\data_path/si_w[13] ), .A1(n732), .B0(n544), .B1(IM_Q[13]), 
        .Y(n390) );
  AO22X1 U792 ( .A0(n725), .A1(\data_path/si_w[14] ), .B0(n724), .B1(
        curr_time[14]), .Y(n325) );
  AOI2BB2X1 U793 ( .B0(n467), .B1(n529), .A0N(n467), .A1N(curr_photo_addr[14]), 
        .Y(n385) );
  AOI2BB2X1 U794 ( .B0(n466), .B1(n529), .A0N(n466), .A1N(fb_addr[14]), .Y(
        n386) );
  AO22X1 U795 ( .A0(\data_path/si_w[14] ), .A1(n732), .B0(n544), .B1(IM_Q[14]), 
        .Y(n387) );
  AO22X1 U796 ( .A0(n725), .A1(\data_path/si_w[15] ), .B0(n724), .B1(
        curr_time[15]), .Y(n324) );
  AOI2BB2X1 U797 ( .B0(n467), .B1(n525), .A0N(n467), .A1N(curr_photo_addr[15]), 
        .Y(n382) );
  AOI2BB2X1 U798 ( .B0(n466), .B1(n525), .A0N(en_fb_addr), .A1N(fb_addr[15]), 
        .Y(n383) );
  AO22X1 U799 ( .A0(\data_path/si_w[15] ), .A1(n732), .B0(n544), .B1(IM_Q[15]), 
        .Y(n384) );
  AOI2BB2X1 U800 ( .B0(n467), .B1(n527), .A0N(n467), .A1N(curr_photo_addr[17]), 
        .Y(n379) );
  AOI2BB2X1 U801 ( .B0(n466), .B1(n527), .A0N(en_fb_addr), .A1N(fb_addr[17]), 
        .Y(n380) );
  AO22X1 U802 ( .A0(\data_path/si_w[17] ), .A1(n732), .B0(n544), .B1(IM_Q[17]), 
        .Y(n381) );
  OAI222XL U803 ( .A0(n730), .A1(n727), .B0(n540), .B1(en_so), .C0(n726), .C1(
        n729), .Y(n348) );
  AOI2BB2X1 U804 ( .B0(n467), .B1(n526), .A0N(n467), .A1N(curr_photo_addr[18]), 
        .Y(n376) );
  AOI2BB2X1 U805 ( .B0(n466), .B1(n526), .A0N(en_fb_addr), .A1N(fb_addr[18]), 
        .Y(n377) );
  AO22X1 U806 ( .A0(\data_path/si_w[18] ), .A1(n732), .B0(n544), .B1(IM_Q[18]), 
        .Y(n378) );
  OAI2BB2XL U807 ( .B0(n730), .B1(n729), .A0N(im_d_w_19), .A1N(n728), .Y(n347)
         );
  AOI2BB2X1 U808 ( .B0(n467), .B1(n528), .A0N(n467), .A1N(curr_photo_addr[19]), 
        .Y(n373) );
  AOI2BB2X1 U809 ( .B0(n466), .B1(n528), .A0N(en_fb_addr), .A1N(fb_addr[19]), 
        .Y(n374) );
  AO22X1 U810 ( .A0(\data_path/si_w[19] ), .A1(n732), .B0(n544), .B1(IM_Q[19]), 
        .Y(n375) );
  AO22X1 U811 ( .A0(\data_path/si_w[20] ), .A1(n732), .B0(n544), .B1(IM_Q[20]), 
        .Y(n372) );
  AO22X1 U812 ( .A0(\data_path/si_w[21] ), .A1(n732), .B0(n544), .B1(IM_Q[21]), 
        .Y(n371) );
  AO22X1 U813 ( .A0(\data_path/si_w[22] ), .A1(n732), .B0(n544), .B1(IM_Q[22]), 
        .Y(n370) );
  AO22X1 U814 ( .A0(\data_path/si_w[23] ), .A1(n732), .B0(n544), .B1(IM_Q[23]), 
        .Y(n369) );
  AO22X1 U815 ( .A0(n467), .A1(\data_path/si_w[16] ), .B0(n547), .B1(
        curr_photo_addr[16]), .Y(n11) );
  AO22X1 U816 ( .A0(en_fb_addr), .A1(\data_path/si_w[16] ), .B0(n548), .B1(
        fb_addr[16]), .Y(n12) );
  AOI2BB2X1 U817 ( .B0(n467), .B1(n501), .A0N(n467), .A1N(curr_photo_addr[8]), 
        .Y(n13) );
  AOI2BB2X1 U818 ( .B0(n466), .B1(n501), .A0N(n466), .A1N(fb_addr[8]), .Y(n14)
         );
  AOI2BB2X1 U819 ( .B0(n467), .B1(n510), .A0N(n467), .A1N(curr_photo_addr[4]), 
        .Y(n15) );
  AOI2BB2X1 U820 ( .B0(n466), .B1(n510), .A0N(en_fb_addr), .A1N(fb_addr[4]), 
        .Y(n16) );
  AOI2BB2X1 U821 ( .B0(n467), .B1(n511), .A0N(n467), .A1N(curr_photo_addr[2]), 
        .Y(n17) );
  AOI2BB2X1 U822 ( .B0(n466), .B1(n511), .A0N(en_fb_addr), .A1N(fb_addr[2]), 
        .Y(n18) );
  AOI2BB2X1 U823 ( .B0(n467), .B1(n505), .A0N(n467), .A1N(curr_photo_addr[1]), 
        .Y(n19) );
  AOI2BB2X1 U824 ( .B0(n466), .B1(n505), .A0N(en_fb_addr), .A1N(fb_addr[1]), 
        .Y(n20) );
  OAI22XL U825 ( .A0(\data_path/si_w[0] ), .A1(n505), .B0(n516), .B1(
        \data_path/si_w[1] ), .Y(n733) );
  OAI21XL U826 ( .A0(en_curr_photo_size), .A1(n537), .B0(n735), .Y(n23) );
endmodule

