
module CONT ( clk, reset, im_wen_n, cr_a, curr_time, fb_addr, photo_num, 
        curr_photo_addr, curr_photo_size, en_si, en_init_time, en_fb_addr, 
        en_photo_num, en_curr_photo_addr, en_curr_photo_size, en_so, si_sel, 
        init_time_mux_sel, sftr_n, so_mux_sel, expand_sel, \im_a[19]_BAR , 
        \im_a[18]_BAR , \im_a[17]_BAR , \im_a[16]_BAR , \im_a[15]_BAR , 
        \im_a[14]_BAR , \im_a[13]_BAR , \im_a[12]_BAR , \im_a[11]_BAR , 
        \im_a[10]_BAR , \im_a[9]_BAR , \im_a[8]_BAR , \im_a[7]_BAR , 
        \im_a[6]_BAR , \im_a[5]_BAR , \im_a[4]_BAR , \im_a[3]_BAR , 
        \im_a[2]_BAR , \im_a[1]_BAR , \im_a[0]_BAR  );
  output [8:0] cr_a;
  input [23:0] curr_time;
  input [19:0] fb_addr;
  input [1:0] photo_num;
  input [19:0] curr_photo_addr;
  input [1:0] curr_photo_size;
  output [1:0] sftr_n;
  output [1:0] so_mux_sel;
  output [3:0] expand_sel;
  input clk, reset;
  output im_wen_n, en_si, en_init_time, en_fb_addr, en_photo_num,
         en_curr_photo_addr, en_curr_photo_size, en_so, si_sel,
         init_time_mux_sel, \im_a[19]_BAR , \im_a[18]_BAR , \im_a[17]_BAR ,
         \im_a[16]_BAR , \im_a[15]_BAR , \im_a[14]_BAR , \im_a[13]_BAR ,
         \im_a[12]_BAR , \im_a[11]_BAR , \im_a[10]_BAR , \im_a[9]_BAR ,
         \im_a[8]_BAR , \im_a[7]_BAR , \im_a[6]_BAR , \im_a[5]_BAR ,
         \im_a[4]_BAR , \im_a[3]_BAR , \im_a[2]_BAR , \im_a[1]_BAR ,
         \im_a[0]_BAR ;
  wire   n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         \next_write_addr_w[0] , \next_cr_y[0] , \h_0[0] , \m_1[3] , \m_0[0] ,
         \s_1[3] , \s_0[0] , N464, N465, N466, N467, N468, N469, N470, N471,
         N472, N473, N474, N475, N476, N477, N478, N479, N480, N481, N579,
         N580, N581, N582, N583, N584, N585, N587, N588, N589, N590, N591,
         N592, N593, N594, N595, N596, N597, N31, N32, N1232, N1233, N1234,
         N1235, N1236, N1237, N1238, N1239, N1446, N1447, N1448, N1449, N1450,
         N1451, N1452, N1453, N1454, N1455, N1456, N1457, N1458, N1459, N1460,
         N1461, N1462, N1463, N1464, N1465, N2061, N2062, N2063, N85,
         next_en_si, N2622, N2644, N2664, N2666, \C163/Z_0 , \C163/Z_1 ,
         \C163/Z_2 , \C163/Z_3 , \C163/Z_4 , \C163/Z_5 , \C163/Z_6 ,
         \C163/Z_7 , \C163/Z_8 , \C163/Z_9 , \C163/Z_10 , \C163/Z_12 ,
         \C163/Z_13 , \C163/Z_15 , \C163/Z_16 , \C163/Z_17 , \C162/DATA3_0 ,
         \C162/DATA3_1 , \C162/DATA3_2 , \C162/DATA3_3 , \C162/DATA3_4 ,
         \C162/DATA3_5 , \C162/DATA3_6 , \C162/DATA3_7 , \C162/DATA3_8 ,
         \C162/DATA3_9 , \C162/DATA3_10 , \C162/DATA3_11 , \C162/DATA3_12 ,
         \C162/DATA3_13 , \C162/DATA3_14 , \C162/DATA3_15 , \C162/DATA3_16 ,
         \C162/DATA3_17 , \C162/DATA3_18 , \C162/DATA3_19 , n14, n28, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n518, n519, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n534, n535, n536,
         n537, \C1/Z_19 , \C1/Z_18 , \C1/Z_17 , \C1/Z_16 , \C1/Z_15 ,
         \C1/Z_14 , \C1/Z_13 , \C1/Z_12 , \C1/Z_11 , \C1/Z_10 , \C1/Z_9 ,
         \C1/Z_8 , \C1/Z_7 , \C1/Z_6 , \C1/Z_5 , \C1/Z_4 ,
         \U3/RSOP_657/C2/Z_19 , \U3/RSOP_657/C2/Z_18 , \U3/RSOP_657/C2/Z_17 ,
         \U3/RSOP_657/C2/Z_16 , \U3/RSOP_657/C2/Z_15 , \U3/RSOP_657/C2/Z_13 ,
         \U3/RSOP_657/C2/Z_12 , \U3/RSOP_657/C2/Z_11 , \U3/RSOP_657/C2/Z_10 ,
         \U3/RSOP_657/C2/Z_9 , \U3/RSOP_657/C2/Z_8 , \U3/RSOP_657/C2/Z_7 ,
         \U3/RSOP_657/C2/Z_6 , \U3/RSOP_657/C2/Z_5 , \U3/RSOP_657/C2/Z_4 ,
         \U3/RSOP_657/C2/Z_3 , \U3/RSOP_657/C2/Z_2 , \U3/RSOP_657/C2/Z_1 ,
         \U3/RSOP_657/C2/Z_0 , \C1/Z_3 , \C1/Z_2 , \C1/Z_1 , \C1/Z_0 ,
         \DP_OP_251J1_126_494/I2 , \DP_OP_251J1_126_494/I3 ,
         \DP_OP_251J1_126_494/n27 , \DP_OP_251J1_126_494/n26 ,
         \DP_OP_251J1_126_494/n25 , \DP_OP_251J1_126_494/n24 ,
         \DP_OP_251J1_126_494/n23 , \DP_OP_251J1_126_494/n21 ,
         \DP_OP_251J1_126_494/n17 , \DP_OP_251J1_126_494/n16 ,
         \DP_OP_251J1_126_494/n8 , \DP_OP_251J1_126_494/n7 ,
         \DP_OP_251J1_126_494/n6 , \DP_OP_251J1_126_494/n5 ,
         \DP_OP_251J1_126_494/n4 , \DP_OP_251J1_126_494/n3 ,
         \DP_OP_251J1_126_494/n2 , \DP_OP_251J1_126_494/n1 ,
         \DP_OP_665J1_134_4923/I2 , \DP_OP_665J1_134_4923/I3 ,
         \DP_OP_665J1_134_4923/I4 , \DP_OP_665J1_134_4923/I7 ,
         \DP_OP_665J1_134_4923/I10 , \DP_OP_665J1_134_4923/n270 ,
         \DP_OP_665J1_134_4923/n269 , \DP_OP_665J1_134_4923/n268 ,
         \DP_OP_665J1_134_4923/n267 , \DP_OP_665J1_134_4923/n266 ,
         \DP_OP_665J1_134_4923/n265 , \DP_OP_665J1_134_4923/n264 ,
         \DP_OP_665J1_134_4923/n263 , \DP_OP_665J1_134_4923/n262 ,
         \DP_OP_665J1_134_4923/n261 , \DP_OP_665J1_134_4923/n260 ,
         \DP_OP_665J1_134_4923/n259 , \DP_OP_665J1_134_4923/n250 ,
         \DP_OP_665J1_134_4923/n249 , \DP_OP_665J1_134_4923/n248 ,
         \DP_OP_665J1_134_4923/n246 , \DP_OP_665J1_134_4923/n245 ,
         \DP_OP_665J1_134_4923/n243 , \DP_OP_665J1_134_4923/n242 ,
         \DP_OP_665J1_134_4923/n241 , \DP_OP_665J1_134_4923/n240 ,
         \DP_OP_665J1_134_4923/n239 , \DP_OP_665J1_134_4923/n238 ,
         \DP_OP_665J1_134_4923/n237 , \DP_OP_665J1_134_4923/n236 ,
         \DP_OP_665J1_134_4923/n235 , \DP_OP_665J1_134_4923/n234 ,
         \DP_OP_665J1_134_4923/n233 , \DP_OP_665J1_134_4923/n232 ,
         \DP_OP_665J1_134_4923/n231 , \DP_OP_665J1_134_4923/n230 ,
         \DP_OP_665J1_134_4923/n229 , \DP_OP_665J1_134_4923/n228 ,
         \DP_OP_665J1_134_4923/n227 , \DP_OP_665J1_134_4923/n226 ,
         \DP_OP_665J1_134_4923/n225 , \DP_OP_665J1_134_4923/n224 ,
         \DP_OP_665J1_134_4923/n223 , \DP_OP_665J1_134_4923/n222 ,
         \DP_OP_665J1_134_4923/n221 , \DP_OP_665J1_134_4923/n220 ,
         \DP_OP_665J1_134_4923/n219 , \DP_OP_665J1_134_4923/n218 ,
         \DP_OP_665J1_134_4923/n217 , \DP_OP_665J1_134_4923/n216 ,
         \DP_OP_665J1_134_4923/n215 , \DP_OP_665J1_134_4923/n214 ,
         \DP_OP_665J1_134_4923/n213 , \DP_OP_665J1_134_4923/n206 ,
         \DP_OP_665J1_134_4923/n205 , \DP_OP_665J1_134_4923/n203 ,
         \DP_OP_665J1_134_4923/n202 , \DP_OP_665J1_134_4923/n200 ,
         \DP_OP_665J1_134_4923/n199 , \DP_OP_665J1_134_4923/n198 ,
         \DP_OP_665J1_134_4923/n197 , \DP_OP_665J1_134_4923/n196 ,
         \DP_OP_665J1_134_4923/n195 , \DP_OP_665J1_134_4923/n194 ,
         \DP_OP_665J1_134_4923/n193 , \DP_OP_665J1_134_4923/n192 ,
         \DP_OP_665J1_134_4923/n190 , \DP_OP_665J1_134_4923/n187 ,
         \DP_OP_665J1_134_4923/n184 , \DP_OP_665J1_134_4923/n183 ,
         \DP_OP_665J1_134_4923/n182 , \DP_OP_665J1_134_4923/n181 ,
         \DP_OP_665J1_134_4923/n180 , \DP_OP_665J1_134_4923/n179 ,
         \DP_OP_665J1_134_4923/n178 , \DP_OP_665J1_134_4923/n177 ,
         \DP_OP_665J1_134_4923/n176 , \DP_OP_665J1_134_4923/n175 ,
         \DP_OP_665J1_134_4923/n173 , \DP_OP_665J1_134_4923/n172 ,
         \DP_OP_665J1_134_4923/n171 , \DP_OP_665J1_134_4923/n170 ,
         \DP_OP_665J1_134_4923/n169 , \DP_OP_665J1_134_4923/n168 ,
         \DP_OP_665J1_134_4923/n167 , \DP_OP_665J1_134_4923/n166 ,
         \DP_OP_665J1_134_4923/n165 , \DP_OP_665J1_134_4923/n164 ,
         \DP_OP_665J1_134_4923/n163 , \DP_OP_665J1_134_4923/n162 ,
         \DP_OP_665J1_134_4923/n161 , \DP_OP_665J1_134_4923/n160 ,
         \DP_OP_665J1_134_4923/n159 , \DP_OP_665J1_134_4923/n158 ,
         \DP_OP_665J1_134_4923/n157 , \DP_OP_665J1_134_4923/n156 ,
         \DP_OP_665J1_134_4923/n155 , \DP_OP_665J1_134_4923/n154 ,
         \DP_OP_665J1_134_4923/n153 , \DP_OP_665J1_134_4923/n152 ,
         \DP_OP_665J1_134_4923/n151 , \DP_OP_665J1_134_4923/n150 ,
         \DP_OP_665J1_134_4923/n149 , \DP_OP_665J1_134_4923/n148 ,
         \DP_OP_665J1_134_4923/n147 , \DP_OP_665J1_134_4923/n146 ,
         \DP_OP_665J1_134_4923/n144 , \DP_OP_665J1_134_4923/n143 ,
         \DP_OP_665J1_134_4923/n142 , \DP_OP_665J1_134_4923/n141 ,
         \DP_OP_665J1_134_4923/n140 , \DP_OP_665J1_134_4923/n139 ,
         \DP_OP_665J1_134_4923/n138 , \DP_OP_665J1_134_4923/n137 ,
         \DP_OP_665J1_134_4923/n136 , \DP_OP_665J1_134_4923/n135 ,
         \DP_OP_665J1_134_4923/n134 , \DP_OP_665J1_134_4923/n133 ,
         \DP_OP_665J1_134_4923/n132 , \DP_OP_665J1_134_4923/n131 ,
         \DP_OP_665J1_134_4923/n130 , \DP_OP_665J1_134_4923/n129 ,
         \DP_OP_665J1_134_4923/n128 , \DP_OP_665J1_134_4923/n127 ,
         \DP_OP_665J1_134_4923/n126 , \DP_OP_665J1_134_4923/n125 ,
         \DP_OP_665J1_134_4923/n124 , \DP_OP_665J1_134_4923/n123 ,
         \DP_OP_665J1_134_4923/n122 , \DP_OP_665J1_134_4923/n121 ,
         \DP_OP_665J1_134_4923/n120 , \DP_OP_665J1_134_4923/n119 ,
         \DP_OP_665J1_134_4923/n118 , \DP_OP_665J1_134_4923/n117 ,
         \DP_OP_665J1_134_4923/n116 , \DP_OP_665J1_134_4923/n115 ,
         \DP_OP_665J1_134_4923/n114 , \DP_OP_665J1_134_4923/n113 ,
         \DP_OP_665J1_134_4923/n112 , \DP_OP_665J1_134_4923/n111 ,
         \DP_OP_665J1_134_4923/n110 , \DP_OP_665J1_134_4923/n105 ,
         \DP_OP_665J1_134_4923/n104 , \DP_OP_665J1_134_4923/n103 ,
         \DP_OP_665J1_134_4923/n102 , \DP_OP_665J1_134_4923/n101 ,
         \DP_OP_665J1_134_4923/n100 , \DP_OP_665J1_134_4923/n99 ,
         \DP_OP_665J1_134_4923/n98 , \DP_OP_665J1_134_4923/n93 ,
         \DP_OP_665J1_134_4923/n92 , \DP_OP_665J1_134_4923/n91 ,
         \DP_OP_665J1_134_4923/n90 , \DP_OP_665J1_134_4923/n89 ,
         \DP_OP_665J1_134_4923/n88 , \DP_OP_665J1_134_4923/n87 ,
         \DP_OP_665J1_134_4923/n86 , \DP_OP_665J1_134_4923/n85 ,
         \DP_OP_665J1_134_4923/n84 , \DP_OP_665J1_134_4923/n83 ,
         \DP_OP_665J1_134_4923/n82 , \DP_OP_665J1_134_4923/n77 ,
         \DP_OP_665J1_134_4923/n76 , \DP_OP_665J1_134_4923/n75 ,
         \DP_OP_665J1_134_4923/n74 , \DP_OP_665J1_134_4923/n73 ,
         \DP_OP_665J1_134_4923/n72 , \DP_OP_665J1_134_4923/n71 ,
         \DP_OP_665J1_134_4923/n70 , \DP_OP_665J1_134_4923/n69 ,
         \DP_OP_665J1_134_4923/n68 , \DP_OP_665J1_134_4923/n67 ,
         \DP_OP_665J1_134_4923/n66 , \DP_OP_665J1_134_4923/n65 ,
         \DP_OP_665J1_134_4923/n64 , \DP_OP_665J1_134_4923/n63 ,
         \DP_OP_665J1_134_4923/n62 , \DP_OP_665J1_134_4923/n61 ,
         \DP_OP_665J1_134_4923/n60 , \DP_OP_665J1_134_4923/n59 ,
         \DP_OP_665J1_134_4923/n58 , \DP_OP_665J1_134_4923/n57 ,
         \DP_OP_665J1_134_4923/n56 , \DP_OP_665J1_134_4923/n55 ,
         \DP_OP_665J1_134_4923/n54 , \DP_OP_665J1_134_4923/n53 ,
         \DP_OP_665J1_134_4923/n52 , \DP_OP_665J1_134_4923/n51 ,
         \DP_OP_665J1_134_4923/n50 , \DP_OP_665J1_134_4923/n49 ,
         \DP_OP_665J1_134_4923/n48 , \DP_OP_665J1_134_4923/n47 ,
         \DP_OP_665J1_134_4923/n46 , \DP_OP_665J1_134_4923/n45 ,
         \DP_OP_665J1_134_4923/n44 , \DP_OP_665J1_134_4923/n43 ,
         \DP_OP_665J1_134_4923/n42 , \DP_OP_665J1_134_4923/n41 ,
         \DP_OP_665J1_134_4923/n40 , \DP_OP_665J1_134_4923/n39 ,
         \DP_OP_665J1_134_4923/n38 , \DP_OP_665J1_134_4923/n37 ,
         \DP_OP_665J1_134_4923/n36 , \DP_OP_665J1_134_4923/n35 ,
         \DP_OP_665J1_134_4923/n34 , \DP_OP_665J1_134_4923/n33 ,
         \DP_OP_665J1_134_4923/n32 , \DP_OP_665J1_134_4923/n31 ,
         \DP_OP_665J1_134_4923/n30 , \DP_OP_665J1_134_4923/n29 ,
         \DP_OP_665J1_134_4923/n28 , \DP_OP_665J1_134_4923/n27 ,
         \DP_OP_665J1_134_4923/n26 , \DP_OP_665J1_134_4923/n25 ,
         \DP_OP_665J1_134_4923/n24 , \DP_OP_665J1_134_4923/n23 ,
         \DP_OP_665J1_134_4923/n22 , \DP_OP_665J1_134_4923/n21 ,
         \DP_OP_665J1_134_4923/n20 , \DP_OP_665J1_134_4923/n19 ,
         \DP_OP_665J1_134_4923/n18 , \DP_OP_665J1_134_4923/n17 ,
         \DP_OP_665J1_134_4923/n16 , \DP_OP_665J1_134_4923/n15 ,
         \DP_OP_665J1_134_4923/n14 , \DP_OP_665J1_134_4923/n13 ,
         \DP_OP_665J1_134_4923/n12 , \DP_OP_665J1_134_4923/n11 ,
         \DP_OP_665J1_134_4923/n10 , \DP_OP_665J1_134_4923/n9 ,
         \DP_OP_665J1_134_4923/n8 , \DP_OP_665J1_134_4923/n7 ,
         \DP_OP_665J1_134_4923/n6 , \DP_OP_665J1_134_4923/n5 ,
         \DP_OP_665J1_134_4923/n4 , \DP_OP_665J1_134_4923/n3 ,
         \DP_OP_665J1_134_4923/n2 , \DP_OP_665J1_134_4923/n1 , \intadd_3/A[4] ,
         \intadd_3/A[3] , \intadd_3/A[2] , \intadd_3/A[1] , \intadd_3/A[0] ,
         \intadd_3/B[6] , \intadd_3/B[5] , \intadd_3/B[4] , \intadd_3/B[3] ,
         \intadd_3/B[2] , \intadd_3/B[1] , \intadd_3/B[0] , \intadd_3/CI ,
         \intadd_3/SUM[6] , \intadd_3/SUM[5] , \intadd_3/SUM[4] ,
         \intadd_3/SUM[3] , \intadd_3/SUM[2] , \intadd_3/SUM[1] ,
         \intadd_3/SUM[0] , \intadd_3/n7 , \intadd_3/n6 , \intadd_3/n5 ,
         \intadd_3/n4 , \intadd_3/n3 , \intadd_3/n2 , \intadd_3/n1 ,
         \intadd_4/A[2] , \intadd_4/A[1] , \intadd_4/B[3] , \intadd_4/B[1] ,
         \intadd_4/SUM[3] , \intadd_4/SUM[2] , \intadd_4/SUM[1] ,
         \intadd_4/SUM[0] , \intadd_4/n4 , \intadd_4/n3 , n1, n2, n3, n4, n5,
         n6, n7, n8, n10, n12, n15, n17, n19, n21, n23, n25, n27, n30, n32,
         n34, n36, n38, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n136, n138, n140, n142, n144, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n219, n221, n222, n223, n224, n225, n226, n227, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n520, n521, n533, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340;
  wire   [2:0] next_state;
  wire   [2:0] state;
  wire   [19:0] work_cntr;
  wire   [19:0] next_work_cntr;
  wire   [19:0] global_cntr;
  wire   [19:0] next_glb_cntr;
  wire   [19:0] write_addr;
  wire   [19:0] write_cntr;
  wire   [8:0] next_cr_x;
  wire   [3:0] h_1;
  wire   [19:0] read_cntr;
  wire   [8:0] cr_read_cntr;
  wire   [1:0] curr_photo;
  wire   [1:0] next_photo;
  assign \h_0[0]  = curr_time[16];
  assign \m_0[0]  = curr_time[8];
  assign \s_0[0]  = curr_time[0];
  assign en_init_time = N2622;
  assign en_curr_photo_addr = N2644;
  assign en_curr_photo_size = N2664;
  assign init_time_mux_sel = N2666;

  DFFSX1 en_si_reg ( .D(next_en_si), .CK(clk), .SN(n275), .Q(en_si) );
  ADDHXL \DP_OP_251J1_126_494/U16  ( .A(\C1/Z_0 ), .B(\C1/Z_1 ), .CO(
        \DP_OP_251J1_126_494/n8 ), .S(\DP_OP_251J1_126_494/n23 ) );
  ADDFXL \DP_OP_251J1_126_494/U15  ( .A(\C1/Z_2 ), .B(\C1/Z_1 ), .CI(
        \DP_OP_251J1_126_494/n8 ), .CO(\DP_OP_251J1_126_494/n7 ), .S(
        \DP_OP_251J1_126_494/n24 ) );
  ADDFXL \DP_OP_251J1_126_494/U14  ( .A(\C1/Z_3 ), .B(\C1/Z_2 ), .CI(
        \DP_OP_251J1_126_494/n7 ), .CO(\DP_OP_251J1_126_494/n6 ), .S(
        \DP_OP_251J1_126_494/n25 ) );
  ADDHXL \DP_OP_251J1_126_494/U13  ( .A(\C1/Z_3 ), .B(\DP_OP_251J1_126_494/n6 ), .CO(\DP_OP_251J1_126_494/n27 ), .S(\DP_OP_251J1_126_494/n26 ) );
  AO21X1 \DP_OP_251J1_126_494/U11  ( .A0(\DP_OP_251J1_126_494/n23 ), .A1(
        \DP_OP_251J1_126_494/I3 ), .B0(\DP_OP_251J1_126_494/I2 ), .Y(
        \DP_OP_251J1_126_494/n17 ) );
  ADDHXL \DP_OP_665J1_134_4923/U245  ( .A(write_addr[11]), .B(
        \DP_OP_665J1_134_4923/n200 ), .CO(\DP_OP_665J1_134_4923/n199 ), .S(
        \DP_OP_665J1_134_4923/n261 ) );
  ADDHXL \DP_OP_665J1_134_4923/U244  ( .A(write_addr[12]), .B(
        \DP_OP_665J1_134_4923/n199 ), .CO(\DP_OP_665J1_134_4923/n198 ), .S(
        \DP_OP_665J1_134_4923/n262 ) );
  ADDHXL \DP_OP_665J1_134_4923/U243  ( .A(write_addr[13]), .B(
        \DP_OP_665J1_134_4923/n198 ), .CO(\DP_OP_665J1_134_4923/n197 ), .S(
        \DP_OP_665J1_134_4923/n263 ) );
  ADDHXL \DP_OP_665J1_134_4923/U242  ( .A(write_addr[14]), .B(
        \DP_OP_665J1_134_4923/n197 ), .CO(\DP_OP_665J1_134_4923/n196 ), .S(
        \DP_OP_665J1_134_4923/n264 ) );
  ADDHXL \DP_OP_665J1_134_4923/U241  ( .A(write_addr[15]), .B(
        \DP_OP_665J1_134_4923/n196 ), .CO(\DP_OP_665J1_134_4923/n195 ), .S(
        \DP_OP_665J1_134_4923/n265 ) );
  ADDHXL \DP_OP_665J1_134_4923/U240  ( .A(write_addr[16]), .B(
        \DP_OP_665J1_134_4923/n195 ), .CO(\DP_OP_665J1_134_4923/n194 ), .S(
        \DP_OP_665J1_134_4923/n266 ) );
  ADDHXL \DP_OP_665J1_134_4923/U239  ( .A(n271), .B(
        \DP_OP_665J1_134_4923/n194 ), .CO(\DP_OP_665J1_134_4923/n193 ), .S(
        \DP_OP_665J1_134_4923/n267 ) );
  ADDHXL \DP_OP_665J1_134_4923/U238  ( .A(write_addr[18]), .B(
        \DP_OP_665J1_134_4923/n193 ), .CO(\DP_OP_665J1_134_4923/n192 ), .S(
        \DP_OP_665J1_134_4923/n268 ) );
  ADDHXL \DP_OP_665J1_134_4923/U237  ( .A(write_addr[19]), .B(
        \DP_OP_665J1_134_4923/n192 ), .CO(\DP_OP_665J1_134_4923/n270 ), .S(
        \DP_OP_665J1_134_4923/n269 ) );
  ADDHXL \DP_OP_665J1_134_4923/U218  ( .A(write_addr[19]), .B(
        \DP_OP_665J1_134_4923/n175 ), .CO(N481), .S(N480) );
  ADDFXL \DP_OP_665J1_134_4923/U204  ( .A(N579), .B(fb_addr[1]), .CI(
        \DP_OP_665J1_134_4923/n164 ), .CO(\DP_OP_665J1_134_4923/n163 ), .S(
        N1447) );
  ADDFXL \DP_OP_665J1_134_4923/U203  ( .A(N580), .B(fb_addr[2]), .CI(
        \DP_OP_665J1_134_4923/n163 ), .CO(\DP_OP_665J1_134_4923/n162 ), .S(
        N1448) );
  ADDFXL \DP_OP_665J1_134_4923/U202  ( .A(N581), .B(fb_addr[3]), .CI(
        \DP_OP_665J1_134_4923/n162 ), .CO(\DP_OP_665J1_134_4923/n161 ), .S(
        N1449) );
  ADDFXL \DP_OP_665J1_134_4923/U201  ( .A(n272), .B(fb_addr[4]), .CI(
        \DP_OP_665J1_134_4923/n161 ), .CO(\DP_OP_665J1_134_4923/n160 ), .S(
        N1450) );
  ADDFXL \DP_OP_665J1_134_4923/U200  ( .A(N583), .B(fb_addr[5]), .CI(
        \DP_OP_665J1_134_4923/n160 ), .CO(\DP_OP_665J1_134_4923/n159 ), .S(
        N1451) );
  ADDFXL \DP_OP_665J1_134_4923/U199  ( .A(N584), .B(fb_addr[6]), .CI(
        \DP_OP_665J1_134_4923/n159 ), .CO(\DP_OP_665J1_134_4923/n158 ), .S(
        N1452) );
  ADDFXL \DP_OP_665J1_134_4923/U198  ( .A(N585), .B(fb_addr[7]), .CI(
        \DP_OP_665J1_134_4923/n158 ), .CO(\DP_OP_665J1_134_4923/n157 ), .S(
        N1453) );
  ADDFXL \DP_OP_665J1_134_4923/U197  ( .A(write_addr[8]), .B(fb_addr[8]), .CI(
        \DP_OP_665J1_134_4923/n157 ), .CO(\DP_OP_665J1_134_4923/n156 ), .S(
        N1454) );
  ADDFXL \DP_OP_665J1_134_4923/U196  ( .A(write_addr[9]), .B(fb_addr[9]), .CI(
        \DP_OP_665J1_134_4923/n156 ), .CO(\DP_OP_665J1_134_4923/n155 ), .S(
        N1455) );
  ADDFXL \DP_OP_665J1_134_4923/U195  ( .A(write_addr[10]), .B(fb_addr[10]), 
        .CI(\DP_OP_665J1_134_4923/n155 ), .CO(\DP_OP_665J1_134_4923/n154 ), 
        .S(N1456) );
  ADDFXL \DP_OP_665J1_134_4923/U194  ( .A(write_addr[11]), .B(fb_addr[11]), 
        .CI(\DP_OP_665J1_134_4923/n154 ), .CO(\DP_OP_665J1_134_4923/n153 ), 
        .S(N1457) );
  ADDFXL \DP_OP_665J1_134_4923/U193  ( .A(write_addr[12]), .B(fb_addr[12]), 
        .CI(\DP_OP_665J1_134_4923/n153 ), .CO(\DP_OP_665J1_134_4923/n152 ), 
        .S(N1458) );
  ADDFXL \DP_OP_665J1_134_4923/U192  ( .A(write_addr[13]), .B(fb_addr[13]), 
        .CI(\DP_OP_665J1_134_4923/n152 ), .CO(\DP_OP_665J1_134_4923/n151 ), 
        .S(N1459) );
  ADDFXL \DP_OP_665J1_134_4923/U191  ( .A(write_addr[14]), .B(fb_addr[14]), 
        .CI(\DP_OP_665J1_134_4923/n151 ), .CO(\DP_OP_665J1_134_4923/n150 ), 
        .S(N1460) );
  ADDFXL \DP_OP_665J1_134_4923/U190  ( .A(write_addr[15]), .B(fb_addr[15]), 
        .CI(\DP_OP_665J1_134_4923/n150 ), .CO(\DP_OP_665J1_134_4923/n149 ), 
        .S(N1461) );
  ADDFXL \DP_OP_665J1_134_4923/U189  ( .A(write_addr[16]), .B(fb_addr[16]), 
        .CI(\DP_OP_665J1_134_4923/n149 ), .CO(\DP_OP_665J1_134_4923/n148 ), 
        .S(N1462) );
  ADDFXL \DP_OP_665J1_134_4923/U188  ( .A(n271), .B(fb_addr[17]), .CI(
        \DP_OP_665J1_134_4923/n148 ), .CO(\DP_OP_665J1_134_4923/n147 ), .S(
        N1463) );
  ADDFXL \DP_OP_665J1_134_4923/U187  ( .A(write_addr[18]), .B(fb_addr[18]), 
        .CI(\DP_OP_665J1_134_4923/n147 ), .CO(\DP_OP_665J1_134_4923/n146 ), 
        .S(N1464) );
  AO22X1 \DP_OP_665J1_134_4923/U22  ( .A0(N1465), .A1(si_sel), .B0(
        \DP_OP_665J1_134_4923/I10 ), .B1(\U3/RSOP_657/C2/Z_19 ), .Y(
        \DP_OP_665J1_134_4923/n232 ) );
  ADDHXL \DP_OP_665J1_134_4923/U21  ( .A(n677), .B(\DP_OP_665J1_134_4923/n213 ), .CO(\DP_OP_665J1_134_4923/n20 ), .S(\C162/DATA3_0 ) );
  ADDFXL \DP_OP_665J1_134_4923/U20  ( .A(\DP_OP_665J1_134_4923/n20 ), .B(n678), 
        .CI(\DP_OP_665J1_134_4923/n214 ), .CO(\DP_OP_665J1_134_4923/n19 ), .S(
        \C162/DATA3_1 ) );
  ADDFXL \DP_OP_665J1_134_4923/U19  ( .A(\DP_OP_665J1_134_4923/n215 ), .B(n679), .CI(\DP_OP_665J1_134_4923/n19 ), .CO(\DP_OP_665J1_134_4923/n18 ), .S(
        \C162/DATA3_2 ) );
  ADDFXL \DP_OP_665J1_134_4923/U18  ( .A(\DP_OP_665J1_134_4923/n216 ), .B(n680), .CI(\DP_OP_665J1_134_4923/n18 ), .CO(\DP_OP_665J1_134_4923/n17 ), .S(
        \C162/DATA3_3 ) );
  ADDFXL \DP_OP_665J1_134_4923/U17  ( .A(\DP_OP_665J1_134_4923/n217 ), .B(
        \C1/Z_4 ), .CI(\DP_OP_665J1_134_4923/n17 ), .CO(
        \DP_OP_665J1_134_4923/n16 ), .S(\C162/DATA3_4 ) );
  ADDFXL \DP_OP_665J1_134_4923/U16  ( .A(\DP_OP_665J1_134_4923/n218 ), .B(
        \C1/Z_5 ), .CI(\DP_OP_665J1_134_4923/n16 ), .CO(
        \DP_OP_665J1_134_4923/n15 ), .S(\C162/DATA3_5 ) );
  ADDFXL \DP_OP_665J1_134_4923/U15  ( .A(\DP_OP_665J1_134_4923/n219 ), .B(
        \C1/Z_6 ), .CI(\DP_OP_665J1_134_4923/n15 ), .CO(
        \DP_OP_665J1_134_4923/n14 ), .S(\C162/DATA3_6 ) );
  ADDFXL \DP_OP_665J1_134_4923/U14  ( .A(\DP_OP_665J1_134_4923/n220 ), .B(
        \C1/Z_7 ), .CI(\DP_OP_665J1_134_4923/n14 ), .CO(
        \DP_OP_665J1_134_4923/n13 ), .S(\C162/DATA3_7 ) );
  ADDFXL \DP_OP_665J1_134_4923/U13  ( .A(\DP_OP_665J1_134_4923/n221 ), .B(
        \C1/Z_8 ), .CI(\DP_OP_665J1_134_4923/n13 ), .CO(
        \DP_OP_665J1_134_4923/n12 ), .S(\C162/DATA3_8 ) );
  ADDFXL \DP_OP_665J1_134_4923/U12  ( .A(\DP_OP_665J1_134_4923/n222 ), .B(
        \C1/Z_9 ), .CI(\DP_OP_665J1_134_4923/n12 ), .CO(
        \DP_OP_665J1_134_4923/n11 ), .S(\C162/DATA3_9 ) );
  ADDFXL \DP_OP_665J1_134_4923/U11  ( .A(\DP_OP_665J1_134_4923/n223 ), .B(
        \C1/Z_10 ), .CI(\DP_OP_665J1_134_4923/n11 ), .CO(
        \DP_OP_665J1_134_4923/n10 ), .S(\C162/DATA3_10 ) );
  ADDFXL \DP_OP_665J1_134_4923/U10  ( .A(\DP_OP_665J1_134_4923/n224 ), .B(
        \C1/Z_11 ), .CI(\DP_OP_665J1_134_4923/n10 ), .CO(
        \DP_OP_665J1_134_4923/n9 ), .S(\C162/DATA3_11 ) );
  ADDFXL \DP_OP_665J1_134_4923/U9  ( .A(\DP_OP_665J1_134_4923/n225 ), .B(
        \C1/Z_12 ), .CI(\DP_OP_665J1_134_4923/n9 ), .CO(
        \DP_OP_665J1_134_4923/n8 ), .S(\C162/DATA3_12 ) );
  ADDFXL \DP_OP_665J1_134_4923/U8  ( .A(\DP_OP_665J1_134_4923/n226 ), .B(
        \C1/Z_13 ), .CI(\DP_OP_665J1_134_4923/n8 ), .CO(
        \DP_OP_665J1_134_4923/n7 ), .S(\C162/DATA3_13 ) );
  ADDFXL \DP_OP_665J1_134_4923/U7  ( .A(\DP_OP_665J1_134_4923/n227 ), .B(
        \C1/Z_14 ), .CI(\DP_OP_665J1_134_4923/n7 ), .CO(
        \DP_OP_665J1_134_4923/n6 ), .S(\C162/DATA3_14 ) );
  ADDFXL \DP_OP_665J1_134_4923/U6  ( .A(\DP_OP_665J1_134_4923/n228 ), .B(
        \C1/Z_15 ), .CI(\DP_OP_665J1_134_4923/n6 ), .CO(
        \DP_OP_665J1_134_4923/n5 ), .S(\C162/DATA3_15 ) );
  ADDFXL \DP_OP_665J1_134_4923/U5  ( .A(\DP_OP_665J1_134_4923/n229 ), .B(
        \C1/Z_16 ), .CI(\DP_OP_665J1_134_4923/n5 ), .CO(
        \DP_OP_665J1_134_4923/n4 ), .S(\C162/DATA3_16 ) );
  ADDFXL \DP_OP_665J1_134_4923/U4  ( .A(\DP_OP_665J1_134_4923/n230 ), .B(
        \C1/Z_17 ), .CI(\DP_OP_665J1_134_4923/n4 ), .CO(
        \DP_OP_665J1_134_4923/n3 ), .S(\C162/DATA3_17 ) );
  ADDFXL \DP_OP_665J1_134_4923/U3  ( .A(\DP_OP_665J1_134_4923/n231 ), .B(
        \C1/Z_18 ), .CI(\DP_OP_665J1_134_4923/n3 ), .CO(
        \DP_OP_665J1_134_4923/n2 ), .S(\C162/DATA3_18 ) );
  ADDFXL \intadd_3/U8  ( .A(\intadd_3/A[0] ), .B(\intadd_3/B[0] ), .CI(
        \intadd_3/CI ), .CO(\intadd_3/n7 ), .S(\intadd_3/SUM[0] ) );
  ADDFXL \intadd_3/U7  ( .A(\intadd_3/A[1] ), .B(\intadd_3/B[1] ), .CI(
        \intadd_3/n7 ), .CO(\intadd_3/n6 ), .S(\intadd_3/SUM[1] ) );
  ADDFXL \intadd_3/U6  ( .A(\intadd_3/A[2] ), .B(\intadd_3/B[2] ), .CI(
        \intadd_3/n6 ), .CO(\intadd_3/n5 ), .S(\intadd_3/SUM[2] ) );
  ADDFXL \intadd_3/U5  ( .A(\intadd_3/A[3] ), .B(\intadd_3/B[3] ), .CI(
        \intadd_3/n5 ), .CO(\intadd_3/n4 ), .S(\intadd_3/SUM[3] ) );
  ADDFXL \intadd_3/U4  ( .A(\intadd_3/A[4] ), .B(\intadd_3/B[4] ), .CI(
        \intadd_3/n4 ), .CO(\intadd_3/n3 ), .S(\intadd_3/SUM[4] ) );
  ADDFXL \intadd_3/U3  ( .A(n207), .B(\intadd_3/B[5] ), .CI(\intadd_3/n3 ), 
        .CO(\intadd_3/n2 ), .S(\intadd_3/SUM[5] ) );
  ADDFXL \intadd_3/U2  ( .A(n206), .B(\intadd_3/B[6] ), .CI(\intadd_3/n2 ), 
        .CO(\intadd_3/n1 ), .S(\intadd_3/SUM[6] ) );
  ADDFXL \intadd_4/U4  ( .A(\intadd_4/A[1] ), .B(\intadd_4/B[1] ), .CI(
        \intadd_4/n4 ), .CO(\intadd_4/n3 ), .S(\intadd_4/SUM[1] ) );
  DFFRX1 \cr_read_cntr_reg/q_reg[1]  ( .D(n498), .CK(clk), .RN(n274), .Q(N1233), .QN(n259) );
  DFFRX1 \cr_read_cntr_reg/q_reg[8]  ( .D(n491), .CK(clk), .RN(n274), .Q(
        cr_read_cntr[8]), .QN(n258) );
  DFFRX1 \cr_read_cntr_reg/q_reg[2]  ( .D(n497), .CK(clk), .RN(n274), .Q(N1234), .QN(n257) );
  DFFRX1 \cr_read_cntr_reg/q_reg[4]  ( .D(n495), .CK(clk), .RN(n274), .Q(
        cr_read_cntr[4]), .QN(n256) );
  DFFRX1 \cr_read_cntr_reg/q_reg[7]  ( .D(n492), .CK(clk), .RN(n274), .QN(n249) );
  DFFRX1 \write_cntr_reg/q_reg[13]  ( .D(n523), .CK(clk), .RN(n275), .Q(
        write_cntr[13]), .QN(n230) );
  DFFRX1 \write_cntr_reg/q_reg[2]  ( .D(n536), .CK(clk), .RN(n274), .Q(
        write_cntr[2]), .QN(n225) );
  DFFRX1 \cr_read_cntr_reg/q_reg[5]  ( .D(n494), .CK(clk), .RN(n274), .Q(
        cr_read_cntr[5]), .QN(n189) );
  DFFRX1 \write_addr_reg/q_reg[0]  ( .D(n490), .CK(clk), .RN(n274), .Q(
        \next_write_addr_w[0] ), .QN(n237) );
  DFFRX1 \write_addr_reg/q_reg[17]  ( .D(n473), .CK(clk), .RN(n274), .Q(
        write_addr[17]), .QN(n231) );
  DFFRX1 \write_addr_reg/q_reg[4]  ( .D(n486), .CK(clk), .RN(n274), .Q(N582), 
        .QN(n239) );
  DFFRX1 \write_cntr_reg/q_reg[3]  ( .D(n531), .CK(clk), .RN(n274), .Q(
        write_cntr[3]), .QN(n208) );
  DFFRX1 \write_cntr_reg/q_reg[0]  ( .D(n532), .CK(clk), .RN(n274), .Q(
        write_cntr[0]), .QN(n185) );
  DFFRX1 \write_cntr_reg/q_reg[1]  ( .D(n537), .CK(clk), .RN(n274), .Q(
        write_cntr[1]), .QN(n224) );
  DFFRX1 \write_cntr_reg/q_reg[14]  ( .D(n522), .CK(clk), .RN(n709), .Q(
        write_cntr[14]), .QN(n229) );
  DFFRX1 \write_cntr_reg/q_reg[5]  ( .D(n530), .CK(clk), .RN(n274), .Q(
        write_cntr[5]), .QN(n210) );
  NAND2X1 \DP_OP_665J1_134_4923/U106  ( .A(n112), .B(\DP_OP_665J1_134_4923/I2 ), .Y(\DP_OP_665J1_134_4923/n83 ) );
  NAND2X1 \DP_OP_665J1_134_4923/U111  ( .A(N479), .B(\DP_OP_665J1_134_4923/I2 ), .Y(\DP_OP_665J1_134_4923/n87 ) );
  NAND2X1 \DP_OP_665J1_134_4923/U116  ( .A(N478), .B(\DP_OP_665J1_134_4923/I2 ), .Y(\DP_OP_665J1_134_4923/n91 ) );
  NAND2X1 \DP_OP_665J1_134_4923/U126  ( .A(N476), .B(\DP_OP_665J1_134_4923/I2 ), .Y(\DP_OP_665J1_134_4923/n99 ) );
  NAND2X1 \DP_OP_665J1_134_4923/U131  ( .A(N475), .B(\DP_OP_665J1_134_4923/I2 ), .Y(\DP_OP_665J1_134_4923/n103 ) );
  NAND2X1 \DP_OP_665J1_134_4923/U146  ( .A(N472), .B(\DP_OP_665J1_134_4923/I2 ), .Y(\DP_OP_665J1_134_4923/n115 ) );
  NAND2X1 \DP_OP_665J1_134_4923/U151  ( .A(N471), .B(\DP_OP_665J1_134_4923/I2 ), .Y(\DP_OP_665J1_134_4923/n119 ) );
  NAND2X1 \DP_OP_665J1_134_4923/U155  ( .A(N470), .B(\DP_OP_665J1_134_4923/I2 ), .Y(\DP_OP_665J1_134_4923/n122 ) );
  NAND2X1 \DP_OP_665J1_134_4923/U160  ( .A(N469), .B(\DP_OP_665J1_134_4923/I2 ), .Y(\DP_OP_665J1_134_4923/n126 ) );
  NAND2X1 \DP_OP_665J1_134_4923/U164  ( .A(N468), .B(\DP_OP_665J1_134_4923/I2 ), .Y(\DP_OP_665J1_134_4923/n129 ) );
  NAND2X1 \DP_OP_665J1_134_4923/U168  ( .A(N467), .B(\DP_OP_665J1_134_4923/I2 ), .Y(\DP_OP_665J1_134_4923/n132 ) );
  NAND2X1 \DP_OP_665J1_134_4923/U172  ( .A(N466), .B(\DP_OP_665J1_134_4923/I2 ), .Y(\DP_OP_665J1_134_4923/n135 ) );
  NAND2X1 \DP_OP_665J1_134_4923/U176  ( .A(N465), .B(\DP_OP_665J1_134_4923/I2 ), .Y(\DP_OP_665J1_134_4923/n138 ) );
  AOI22X1 \DP_OP_665J1_134_4923/U183  ( .A0(n238), .A1(
        \DP_OP_665J1_134_4923/I3 ), .B0(n238), .B1(\DP_OP_665J1_134_4923/I2 ), 
        .Y(\DP_OP_665J1_134_4923/n143 ) );
  NAND2X1 \DP_OP_665J1_134_4923/U180  ( .A(N464), .B(\DP_OP_665J1_134_4923/I2 ), .Y(\DP_OP_665J1_134_4923/n141 ) );
  ADDHXL \DP_OP_251J1_126_494/U6  ( .A(N31), .B(\DP_OP_251J1_126_494/n16 ), 
        .CO(\DP_OP_251J1_126_494/n5 ), .S(N1235) );
  NAND2XL \DP_OP_665J1_134_4923/U24  ( .A(N1464), .B(si_sel), .Y(
        \DP_OP_665J1_134_4923/n21 ) );
  NAND2XL \DP_OP_665J1_134_4923/U26  ( .A(\DP_OP_665J1_134_4923/I10 ), .B(
        \U3/RSOP_657/C2/Z_18 ), .Y(\DP_OP_665J1_134_4923/n23 ) );
  NAND3XL \DP_OP_665J1_134_4923/U23  ( .A(\DP_OP_665J1_134_4923/n21 ), .B(
        \DP_OP_665J1_134_4923/n22 ), .C(\DP_OP_665J1_134_4923/n23 ), .Y(
        \DP_OP_665J1_134_4923/n231 ) );
  NAND2XL \DP_OP_665J1_134_4923/U28  ( .A(N1463), .B(si_sel), .Y(
        \DP_OP_665J1_134_4923/n24 ) );
  NAND2XL \DP_OP_665J1_134_4923/U105  ( .A(\DP_OP_665J1_134_4923/n269 ), .B(
        \DP_OP_665J1_134_4923/I3 ), .Y(\DP_OP_665J1_134_4923/n82 ) );
  NAND2XL \DP_OP_665J1_134_4923/U107  ( .A(N596), .B(\DP_OP_665J1_134_4923/I4 ), .Y(\DP_OP_665J1_134_4923/n84 ) );
  NAND2XL \DP_OP_665J1_134_4923/U108  ( .A(n106), .B(\C163/Z_17 ), .Y(
        \DP_OP_665J1_134_4923/n85 ) );
  NAND4XL \DP_OP_665J1_134_4923/U104  ( .A(\DP_OP_665J1_134_4923/n82 ), .B(
        \DP_OP_665J1_134_4923/n83 ), .C(\DP_OP_665J1_134_4923/n84 ), .D(
        \DP_OP_665J1_134_4923/n85 ), .Y(\DP_OP_665J1_134_4923/n250 ) );
  NAND2XL \DP_OP_665J1_134_4923/U29  ( .A(\DP_OP_665J1_134_4923/n250 ), .B(
        \DP_OP_665J1_134_4923/I7 ), .Y(\DP_OP_665J1_134_4923/n25 ) );
  NAND2XL \DP_OP_665J1_134_4923/U30  ( .A(\DP_OP_665J1_134_4923/I10 ), .B(
        \U3/RSOP_657/C2/Z_17 ), .Y(\DP_OP_665J1_134_4923/n26 ) );
  NAND3XL \DP_OP_665J1_134_4923/U27  ( .A(\DP_OP_665J1_134_4923/n24 ), .B(
        \DP_OP_665J1_134_4923/n25 ), .C(\DP_OP_665J1_134_4923/n26 ), .Y(
        \DP_OP_665J1_134_4923/n230 ) );
  NAND2XL \DP_OP_665J1_134_4923/U32  ( .A(N1462), .B(si_sel), .Y(
        \DP_OP_665J1_134_4923/n27 ) );
  NAND2XL \DP_OP_665J1_134_4923/U110  ( .A(\DP_OP_665J1_134_4923/n268 ), .B(
        \DP_OP_665J1_134_4923/I3 ), .Y(\DP_OP_665J1_134_4923/n86 ) );
  NAND2XL \DP_OP_665J1_134_4923/U112  ( .A(N595), .B(\DP_OP_665J1_134_4923/I4 ), .Y(\DP_OP_665J1_134_4923/n88 ) );
  NAND2XL \DP_OP_665J1_134_4923/U113  ( .A(n106), .B(\C163/Z_16 ), .Y(
        \DP_OP_665J1_134_4923/n89 ) );
  NAND4XL \DP_OP_665J1_134_4923/U109  ( .A(\DP_OP_665J1_134_4923/n86 ), .B(
        \DP_OP_665J1_134_4923/n87 ), .C(\DP_OP_665J1_134_4923/n88 ), .D(
        \DP_OP_665J1_134_4923/n89 ), .Y(\DP_OP_665J1_134_4923/n249 ) );
  NAND2XL \DP_OP_665J1_134_4923/U33  ( .A(\DP_OP_665J1_134_4923/n249 ), .B(
        \DP_OP_665J1_134_4923/I7 ), .Y(\DP_OP_665J1_134_4923/n28 ) );
  NAND2XL \DP_OP_665J1_134_4923/U34  ( .A(\DP_OP_665J1_134_4923/I10 ), .B(
        \U3/RSOP_657/C2/Z_16 ), .Y(\DP_OP_665J1_134_4923/n29 ) );
  NAND3XL \DP_OP_665J1_134_4923/U31  ( .A(\DP_OP_665J1_134_4923/n27 ), .B(
        \DP_OP_665J1_134_4923/n28 ), .C(\DP_OP_665J1_134_4923/n29 ), .Y(
        \DP_OP_665J1_134_4923/n229 ) );
  NAND2XL \DP_OP_665J1_134_4923/U36  ( .A(N1461), .B(si_sel), .Y(
        \DP_OP_665J1_134_4923/n30 ) );
  NAND2XL \DP_OP_665J1_134_4923/U115  ( .A(\DP_OP_665J1_134_4923/n267 ), .B(
        \DP_OP_665J1_134_4923/I3 ), .Y(\DP_OP_665J1_134_4923/n90 ) );
  NAND2XL \DP_OP_665J1_134_4923/U117  ( .A(N594), .B(\DP_OP_665J1_134_4923/I4 ), .Y(\DP_OP_665J1_134_4923/n92 ) );
  NAND2XL \DP_OP_665J1_134_4923/U118  ( .A(n106), .B(\C163/Z_15 ), .Y(
        \DP_OP_665J1_134_4923/n93 ) );
  NAND4XL \DP_OP_665J1_134_4923/U114  ( .A(\DP_OP_665J1_134_4923/n90 ), .B(
        \DP_OP_665J1_134_4923/n91 ), .C(\DP_OP_665J1_134_4923/n92 ), .D(
        \DP_OP_665J1_134_4923/n93 ), .Y(\DP_OP_665J1_134_4923/n248 ) );
  NAND2XL \DP_OP_665J1_134_4923/U37  ( .A(\DP_OP_665J1_134_4923/n248 ), .B(
        \DP_OP_665J1_134_4923/I7 ), .Y(\DP_OP_665J1_134_4923/n31 ) );
  NAND2XL \DP_OP_665J1_134_4923/U38  ( .A(\DP_OP_665J1_134_4923/I10 ), .B(
        \U3/RSOP_657/C2/Z_15 ), .Y(\DP_OP_665J1_134_4923/n32 ) );
  NAND3XL \DP_OP_665J1_134_4923/U35  ( .A(\DP_OP_665J1_134_4923/n30 ), .B(
        \DP_OP_665J1_134_4923/n31 ), .C(\DP_OP_665J1_134_4923/n32 ), .Y(
        \DP_OP_665J1_134_4923/n228 ) );
  NAND2XL \DP_OP_665J1_134_4923/U40  ( .A(N1460), .B(si_sel), .Y(
        \DP_OP_665J1_134_4923/n33 ) );
  NAND3XL \DP_OP_665J1_134_4923/U39  ( .A(\DP_OP_665J1_134_4923/n33 ), .B(
        \DP_OP_665J1_134_4923/n34 ), .C(\DP_OP_665J1_134_4923/n35 ), .Y(
        \DP_OP_665J1_134_4923/n227 ) );
  NAND2XL \DP_OP_665J1_134_4923/U44  ( .A(N1459), .B(si_sel), .Y(
        \DP_OP_665J1_134_4923/n36 ) );
  NAND2XL \DP_OP_665J1_134_4923/U125  ( .A(\DP_OP_665J1_134_4923/n265 ), .B(
        \DP_OP_665J1_134_4923/I3 ), .Y(\DP_OP_665J1_134_4923/n98 ) );
  NAND2XL \DP_OP_665J1_134_4923/U127  ( .A(N592), .B(\DP_OP_665J1_134_4923/I4 ), .Y(\DP_OP_665J1_134_4923/n100 ) );
  NAND2XL \DP_OP_665J1_134_4923/U128  ( .A(n106), .B(\C163/Z_13 ), .Y(
        \DP_OP_665J1_134_4923/n101 ) );
  NAND4XL \DP_OP_665J1_134_4923/U124  ( .A(\DP_OP_665J1_134_4923/n98 ), .B(
        \DP_OP_665J1_134_4923/n99 ), .C(\DP_OP_665J1_134_4923/n100 ), .D(
        \DP_OP_665J1_134_4923/n101 ), .Y(\DP_OP_665J1_134_4923/n246 ) );
  NAND2XL \DP_OP_665J1_134_4923/U45  ( .A(\DP_OP_665J1_134_4923/n246 ), .B(
        \DP_OP_665J1_134_4923/I7 ), .Y(\DP_OP_665J1_134_4923/n37 ) );
  NAND2XL \DP_OP_665J1_134_4923/U46  ( .A(\DP_OP_665J1_134_4923/I10 ), .B(
        \U3/RSOP_657/C2/Z_13 ), .Y(\DP_OP_665J1_134_4923/n38 ) );
  NAND3XL \DP_OP_665J1_134_4923/U43  ( .A(\DP_OP_665J1_134_4923/n36 ), .B(
        \DP_OP_665J1_134_4923/n37 ), .C(\DP_OP_665J1_134_4923/n38 ), .Y(
        \DP_OP_665J1_134_4923/n226 ) );
  NAND2XL \DP_OP_665J1_134_4923/U48  ( .A(N1458), .B(si_sel), .Y(
        \DP_OP_665J1_134_4923/n39 ) );
  NAND2XL \DP_OP_665J1_134_4923/U130  ( .A(\DP_OP_665J1_134_4923/n264 ), .B(
        \DP_OP_665J1_134_4923/I3 ), .Y(\DP_OP_665J1_134_4923/n102 ) );
  NAND2XL \DP_OP_665J1_134_4923/U132  ( .A(N591), .B(\DP_OP_665J1_134_4923/I4 ), .Y(\DP_OP_665J1_134_4923/n104 ) );
  NAND2XL \DP_OP_665J1_134_4923/U133  ( .A(n106), .B(\C163/Z_12 ), .Y(
        \DP_OP_665J1_134_4923/n105 ) );
  NAND4XL \DP_OP_665J1_134_4923/U129  ( .A(\DP_OP_665J1_134_4923/n102 ), .B(
        \DP_OP_665J1_134_4923/n103 ), .C(\DP_OP_665J1_134_4923/n104 ), .D(
        \DP_OP_665J1_134_4923/n105 ), .Y(\DP_OP_665J1_134_4923/n245 ) );
  NAND2XL \DP_OP_665J1_134_4923/U49  ( .A(\DP_OP_665J1_134_4923/n245 ), .B(
        \DP_OP_665J1_134_4923/I7 ), .Y(\DP_OP_665J1_134_4923/n40 ) );
  NAND2XL \DP_OP_665J1_134_4923/U50  ( .A(\DP_OP_665J1_134_4923/I10 ), .B(
        \U3/RSOP_657/C2/Z_12 ), .Y(\DP_OP_665J1_134_4923/n41 ) );
  NAND3XL \DP_OP_665J1_134_4923/U47  ( .A(\DP_OP_665J1_134_4923/n39 ), .B(
        \DP_OP_665J1_134_4923/n40 ), .C(\DP_OP_665J1_134_4923/n41 ), .Y(
        \DP_OP_665J1_134_4923/n225 ) );
  NAND2XL \DP_OP_665J1_134_4923/U52  ( .A(N1457), .B(si_sel), .Y(
        \DP_OP_665J1_134_4923/n42 ) );
  NAND2XL \DP_OP_665J1_134_4923/U54  ( .A(\DP_OP_665J1_134_4923/I10 ), .B(
        \U3/RSOP_657/C2/Z_11 ), .Y(\DP_OP_665J1_134_4923/n44 ) );
  NAND3XL \DP_OP_665J1_134_4923/U51  ( .A(\DP_OP_665J1_134_4923/n42 ), .B(
        \DP_OP_665J1_134_4923/n43 ), .C(\DP_OP_665J1_134_4923/n44 ), .Y(
        \DP_OP_665J1_134_4923/n224 ) );
  NAND2XL \DP_OP_665J1_134_4923/U56  ( .A(N1456), .B(si_sel), .Y(
        \DP_OP_665J1_134_4923/n45 ) );
  NAND2XL \DP_OP_665J1_134_4923/U140  ( .A(\DP_OP_665J1_134_4923/n262 ), .B(
        \DP_OP_665J1_134_4923/I3 ), .Y(\DP_OP_665J1_134_4923/n110 ) );
  NAND2XL \DP_OP_665J1_134_4923/U142  ( .A(N589), .B(\DP_OP_665J1_134_4923/I4 ), .Y(\DP_OP_665J1_134_4923/n112 ) );
  NAND2XL \DP_OP_665J1_134_4923/U143  ( .A(n106), .B(\C163/Z_10 ), .Y(
        \DP_OP_665J1_134_4923/n113 ) );
  NAND4XL \DP_OP_665J1_134_4923/U139  ( .A(\DP_OP_665J1_134_4923/n110 ), .B(
        \DP_OP_665J1_134_4923/n111 ), .C(\DP_OP_665J1_134_4923/n112 ), .D(
        \DP_OP_665J1_134_4923/n113 ), .Y(\DP_OP_665J1_134_4923/n243 ) );
  NAND2XL \DP_OP_665J1_134_4923/U57  ( .A(\DP_OP_665J1_134_4923/n243 ), .B(
        \DP_OP_665J1_134_4923/I7 ), .Y(\DP_OP_665J1_134_4923/n46 ) );
  NAND2XL \DP_OP_665J1_134_4923/U58  ( .A(\DP_OP_665J1_134_4923/I10 ), .B(
        \U3/RSOP_657/C2/Z_10 ), .Y(\DP_OP_665J1_134_4923/n47 ) );
  NAND3XL \DP_OP_665J1_134_4923/U55  ( .A(\DP_OP_665J1_134_4923/n45 ), .B(
        \DP_OP_665J1_134_4923/n46 ), .C(\DP_OP_665J1_134_4923/n47 ), .Y(
        \DP_OP_665J1_134_4923/n223 ) );
  NAND2XL \DP_OP_665J1_134_4923/U60  ( .A(N1455), .B(si_sel), .Y(
        \DP_OP_665J1_134_4923/n48 ) );
  NAND2XL \DP_OP_665J1_134_4923/U145  ( .A(\DP_OP_665J1_134_4923/n261 ), .B(
        \DP_OP_665J1_134_4923/I3 ), .Y(\DP_OP_665J1_134_4923/n114 ) );
  NAND2XL \DP_OP_665J1_134_4923/U147  ( .A(N588), .B(\DP_OP_665J1_134_4923/I4 ), .Y(\DP_OP_665J1_134_4923/n116 ) );
  NAND2XL \DP_OP_665J1_134_4923/U148  ( .A(n106), .B(\C163/Z_9 ), .Y(
        \DP_OP_665J1_134_4923/n117 ) );
  NAND4XL \DP_OP_665J1_134_4923/U144  ( .A(\DP_OP_665J1_134_4923/n114 ), .B(
        \DP_OP_665J1_134_4923/n115 ), .C(\DP_OP_665J1_134_4923/n116 ), .D(
        \DP_OP_665J1_134_4923/n117 ), .Y(\DP_OP_665J1_134_4923/n242 ) );
  NAND2XL \DP_OP_665J1_134_4923/U61  ( .A(\DP_OP_665J1_134_4923/n242 ), .B(
        \DP_OP_665J1_134_4923/I7 ), .Y(\DP_OP_665J1_134_4923/n49 ) );
  NAND2XL \DP_OP_665J1_134_4923/U62  ( .A(\DP_OP_665J1_134_4923/I10 ), .B(
        \U3/RSOP_657/C2/Z_9 ), .Y(\DP_OP_665J1_134_4923/n50 ) );
  NAND3XL \DP_OP_665J1_134_4923/U59  ( .A(\DP_OP_665J1_134_4923/n48 ), .B(
        \DP_OP_665J1_134_4923/n49 ), .C(\DP_OP_665J1_134_4923/n50 ), .Y(
        \DP_OP_665J1_134_4923/n222 ) );
  NAND2XL \DP_OP_665J1_134_4923/U64  ( .A(N1454), .B(si_sel), .Y(
        \DP_OP_665J1_134_4923/n51 ) );
  NAND2XL \DP_OP_665J1_134_4923/U150  ( .A(\DP_OP_665J1_134_4923/n260 ), .B(
        \DP_OP_665J1_134_4923/I3 ), .Y(\DP_OP_665J1_134_4923/n118 ) );
  NAND2XL \DP_OP_665J1_134_4923/U152  ( .A(N587), .B(\DP_OP_665J1_134_4923/I4 ), .Y(\DP_OP_665J1_134_4923/n120 ) );
  NAND2XL \DP_OP_665J1_134_4923/U153  ( .A(n106), .B(\C163/Z_8 ), .Y(
        \DP_OP_665J1_134_4923/n121 ) );
  NAND4XL \DP_OP_665J1_134_4923/U149  ( .A(\DP_OP_665J1_134_4923/n118 ), .B(
        \DP_OP_665J1_134_4923/n119 ), .C(\DP_OP_665J1_134_4923/n120 ), .D(
        \DP_OP_665J1_134_4923/n121 ), .Y(\DP_OP_665J1_134_4923/n241 ) );
  NAND2XL \DP_OP_665J1_134_4923/U65  ( .A(\DP_OP_665J1_134_4923/n241 ), .B(
        \DP_OP_665J1_134_4923/I7 ), .Y(\DP_OP_665J1_134_4923/n52 ) );
  NAND2XL \DP_OP_665J1_134_4923/U66  ( .A(\DP_OP_665J1_134_4923/I10 ), .B(
        \U3/RSOP_657/C2/Z_8 ), .Y(\DP_OP_665J1_134_4923/n53 ) );
  NAND3XL \DP_OP_665J1_134_4923/U63  ( .A(\DP_OP_665J1_134_4923/n51 ), .B(
        \DP_OP_665J1_134_4923/n52 ), .C(\DP_OP_665J1_134_4923/n53 ), .Y(
        \DP_OP_665J1_134_4923/n221 ) );
  NAND2XL \DP_OP_665J1_134_4923/U68  ( .A(N1453), .B(si_sel), .Y(
        \DP_OP_665J1_134_4923/n54 ) );
  XNOR2XL \DP_OP_665J1_134_4923/U247  ( .A(\DP_OP_665J1_134_4923/n202 ), .B(
        write_addr[9]), .Y(\DP_OP_665J1_134_4923/n259 ) );
  NAND2XL \DP_OP_665J1_134_4923/U156  ( .A(\DP_OP_665J1_134_4923/n259 ), .B(
        \DP_OP_665J1_134_4923/I3 ), .Y(\DP_OP_665J1_134_4923/n123 ) );
  AOI22XL \DP_OP_665J1_134_4923/U157  ( .A0(n244), .A1(
        \DP_OP_665J1_134_4923/I4 ), .B0(n106), .B1(\C163/Z_7 ), .Y(
        \DP_OP_665J1_134_4923/n124 ) );
  NAND3XL \DP_OP_665J1_134_4923/U154  ( .A(\DP_OP_665J1_134_4923/n122 ), .B(
        \DP_OP_665J1_134_4923/n123 ), .C(\DP_OP_665J1_134_4923/n124 ), .Y(
        \DP_OP_665J1_134_4923/n240 ) );
  NAND2XL \DP_OP_665J1_134_4923/U69  ( .A(\DP_OP_665J1_134_4923/n240 ), .B(
        \DP_OP_665J1_134_4923/I7 ), .Y(\DP_OP_665J1_134_4923/n55 ) );
  NAND2XL \DP_OP_665J1_134_4923/U70  ( .A(\DP_OP_665J1_134_4923/I10 ), .B(
        \U3/RSOP_657/C2/Z_7 ), .Y(\DP_OP_665J1_134_4923/n56 ) );
  NAND3XL \DP_OP_665J1_134_4923/U67  ( .A(\DP_OP_665J1_134_4923/n54 ), .B(
        \DP_OP_665J1_134_4923/n55 ), .C(\DP_OP_665J1_134_4923/n56 ), .Y(
        \DP_OP_665J1_134_4923/n220 ) );
  NAND2XL \DP_OP_665J1_134_4923/U72  ( .A(N1452), .B(si_sel), .Y(
        \DP_OP_665J1_134_4923/n57 ) );
  NAND2XL \DP_OP_665J1_134_4923/U159  ( .A(N469), .B(\DP_OP_665J1_134_4923/I3 ), .Y(\DP_OP_665J1_134_4923/n125 ) );
  AOI22XL \DP_OP_665J1_134_4923/U161  ( .A0(n106), .A1(\C163/Z_6 ), .B0(
        \DP_OP_665J1_134_4923/I4 ), .B1(N585), .Y(\DP_OP_665J1_134_4923/n127 )
         );
  NAND3XL \DP_OP_665J1_134_4923/U158  ( .A(\DP_OP_665J1_134_4923/n126 ), .B(
        \DP_OP_665J1_134_4923/n125 ), .C(\DP_OP_665J1_134_4923/n127 ), .Y(
        \DP_OP_665J1_134_4923/n239 ) );
  NAND2XL \DP_OP_665J1_134_4923/U73  ( .A(\DP_OP_665J1_134_4923/n239 ), .B(
        \DP_OP_665J1_134_4923/I7 ), .Y(\DP_OP_665J1_134_4923/n58 ) );
  NAND2XL \DP_OP_665J1_134_4923/U74  ( .A(\DP_OP_665J1_134_4923/I10 ), .B(
        \U3/RSOP_657/C2/Z_6 ), .Y(\DP_OP_665J1_134_4923/n59 ) );
  NAND3XL \DP_OP_665J1_134_4923/U71  ( .A(\DP_OP_665J1_134_4923/n57 ), .B(
        \DP_OP_665J1_134_4923/n58 ), .C(\DP_OP_665J1_134_4923/n59 ), .Y(
        \DP_OP_665J1_134_4923/n219 ) );
  NAND2XL \DP_OP_665J1_134_4923/U76  ( .A(N1451), .B(si_sel), .Y(
        \DP_OP_665J1_134_4923/n60 ) );
  NAND2XL \DP_OP_665J1_134_4923/U163  ( .A(N468), .B(\DP_OP_665J1_134_4923/I3 ), .Y(\DP_OP_665J1_134_4923/n128 ) );
  AOI22XL \DP_OP_665J1_134_4923/U165  ( .A0(n106), .A1(\C163/Z_5 ), .B0(
        \DP_OP_665J1_134_4923/I4 ), .B1(N584), .Y(\DP_OP_665J1_134_4923/n130 )
         );
  NAND3XL \DP_OP_665J1_134_4923/U162  ( .A(\DP_OP_665J1_134_4923/n129 ), .B(
        \DP_OP_665J1_134_4923/n128 ), .C(\DP_OP_665J1_134_4923/n130 ), .Y(
        \DP_OP_665J1_134_4923/n238 ) );
  NAND2XL \DP_OP_665J1_134_4923/U77  ( .A(\DP_OP_665J1_134_4923/n238 ), .B(
        \DP_OP_665J1_134_4923/I7 ), .Y(\DP_OP_665J1_134_4923/n61 ) );
  NAND2XL \DP_OP_665J1_134_4923/U78  ( .A(\DP_OP_665J1_134_4923/I10 ), .B(
        \U3/RSOP_657/C2/Z_5 ), .Y(\DP_OP_665J1_134_4923/n62 ) );
  NAND3XL \DP_OP_665J1_134_4923/U75  ( .A(\DP_OP_665J1_134_4923/n60 ), .B(
        \DP_OP_665J1_134_4923/n61 ), .C(\DP_OP_665J1_134_4923/n62 ), .Y(
        \DP_OP_665J1_134_4923/n218 ) );
  NAND2XL \DP_OP_665J1_134_4923/U80  ( .A(N1450), .B(si_sel), .Y(
        \DP_OP_665J1_134_4923/n63 ) );
  NAND2XL \DP_OP_665J1_134_4923/U167  ( .A(N467), .B(\DP_OP_665J1_134_4923/I3 ), .Y(\DP_OP_665J1_134_4923/n131 ) );
  AOI22XL \DP_OP_665J1_134_4923/U169  ( .A0(n106), .A1(\C163/Z_4 ), .B0(
        \DP_OP_665J1_134_4923/I4 ), .B1(N583), .Y(\DP_OP_665J1_134_4923/n133 )
         );
  NAND3XL \DP_OP_665J1_134_4923/U166  ( .A(\DP_OP_665J1_134_4923/n132 ), .B(
        \DP_OP_665J1_134_4923/n131 ), .C(\DP_OP_665J1_134_4923/n133 ), .Y(
        \DP_OP_665J1_134_4923/n237 ) );
  NAND2XL \DP_OP_665J1_134_4923/U81  ( .A(\DP_OP_665J1_134_4923/n237 ), .B(
        \DP_OP_665J1_134_4923/I7 ), .Y(\DP_OP_665J1_134_4923/n64 ) );
  NAND2XL \DP_OP_665J1_134_4923/U82  ( .A(\DP_OP_665J1_134_4923/I10 ), .B(
        \U3/RSOP_657/C2/Z_4 ), .Y(\DP_OP_665J1_134_4923/n65 ) );
  NAND3XL \DP_OP_665J1_134_4923/U79  ( .A(\DP_OP_665J1_134_4923/n63 ), .B(
        \DP_OP_665J1_134_4923/n64 ), .C(\DP_OP_665J1_134_4923/n65 ), .Y(
        \DP_OP_665J1_134_4923/n217 ) );
  NAND2XL \DP_OP_665J1_134_4923/U84  ( .A(N1449), .B(si_sel), .Y(
        \DP_OP_665J1_134_4923/n66 ) );
  NAND2XL \DP_OP_665J1_134_4923/U171  ( .A(N466), .B(\DP_OP_665J1_134_4923/I3 ), .Y(\DP_OP_665J1_134_4923/n134 ) );
  AOI22XL \DP_OP_665J1_134_4923/U173  ( .A0(n106), .A1(\C163/Z_3 ), .B0(
        \DP_OP_665J1_134_4923/I4 ), .B1(n272), .Y(\DP_OP_665J1_134_4923/n136 )
         );
  NAND3XL \DP_OP_665J1_134_4923/U170  ( .A(\DP_OP_665J1_134_4923/n135 ), .B(
        \DP_OP_665J1_134_4923/n134 ), .C(\DP_OP_665J1_134_4923/n136 ), .Y(
        \DP_OP_665J1_134_4923/n236 ) );
  NAND2XL \DP_OP_665J1_134_4923/U85  ( .A(\DP_OP_665J1_134_4923/n236 ), .B(
        \DP_OP_665J1_134_4923/I7 ), .Y(\DP_OP_665J1_134_4923/n67 ) );
  NAND2XL \DP_OP_665J1_134_4923/U86  ( .A(\DP_OP_665J1_134_4923/I10 ), .B(
        \U3/RSOP_657/C2/Z_3 ), .Y(\DP_OP_665J1_134_4923/n68 ) );
  NAND3XL \DP_OP_665J1_134_4923/U83  ( .A(\DP_OP_665J1_134_4923/n66 ), .B(
        \DP_OP_665J1_134_4923/n67 ), .C(\DP_OP_665J1_134_4923/n68 ), .Y(
        \DP_OP_665J1_134_4923/n216 ) );
  NAND2XL \DP_OP_665J1_134_4923/U88  ( .A(N1448), .B(si_sel), .Y(
        \DP_OP_665J1_134_4923/n69 ) );
  NAND2XL \DP_OP_665J1_134_4923/U175  ( .A(N465), .B(\DP_OP_665J1_134_4923/I3 ), .Y(\DP_OP_665J1_134_4923/n137 ) );
  AOI22XL \DP_OP_665J1_134_4923/U177  ( .A0(n106), .A1(\C163/Z_2 ), .B0(
        \DP_OP_665J1_134_4923/I4 ), .B1(N581), .Y(\DP_OP_665J1_134_4923/n139 )
         );
  NAND3XL \DP_OP_665J1_134_4923/U174  ( .A(\DP_OP_665J1_134_4923/n138 ), .B(
        \DP_OP_665J1_134_4923/n137 ), .C(\DP_OP_665J1_134_4923/n139 ), .Y(
        \DP_OP_665J1_134_4923/n235 ) );
  NAND2XL \DP_OP_665J1_134_4923/U89  ( .A(\DP_OP_665J1_134_4923/n235 ), .B(
        \DP_OP_665J1_134_4923/I7 ), .Y(\DP_OP_665J1_134_4923/n70 ) );
  NAND2XL \DP_OP_665J1_134_4923/U90  ( .A(\DP_OP_665J1_134_4923/I10 ), .B(
        \U3/RSOP_657/C2/Z_2 ), .Y(\DP_OP_665J1_134_4923/n71 ) );
  NAND3XL \DP_OP_665J1_134_4923/U87  ( .A(\DP_OP_665J1_134_4923/n69 ), .B(
        \DP_OP_665J1_134_4923/n70 ), .C(\DP_OP_665J1_134_4923/n71 ), .Y(
        \DP_OP_665J1_134_4923/n215 ) );
  AOI22XL \DP_OP_665J1_134_4923/U184  ( .A0(n106), .A1(\C163/Z_0 ), .B0(
        \DP_OP_665J1_134_4923/I4 ), .B1(N579), .Y(\DP_OP_665J1_134_4923/n144 )
         );
  NAND2XL \DP_OP_665J1_134_4923/U182  ( .A(\DP_OP_665J1_134_4923/n143 ), .B(
        \DP_OP_665J1_134_4923/n144 ), .Y(\DP_OP_665J1_134_4923/n233 ) );
  NAND2XL \DP_OP_665J1_134_4923/U96  ( .A(\DP_OP_665J1_134_4923/n233 ), .B(
        \DP_OP_665J1_134_4923/I7 ), .Y(\DP_OP_665J1_134_4923/n75 ) );
  NAND2XL \DP_OP_665J1_134_4923/U97  ( .A(N1446), .B(si_sel), .Y(
        \DP_OP_665J1_134_4923/n76 ) );
  NAND2XL \DP_OP_665J1_134_4923/U98  ( .A(\DP_OP_665J1_134_4923/I10 ), .B(
        \U3/RSOP_657/C2/Z_0 ), .Y(\DP_OP_665J1_134_4923/n77 ) );
  NAND3XL \DP_OP_665J1_134_4923/U95  ( .A(\DP_OP_665J1_134_4923/n75 ), .B(
        \DP_OP_665J1_134_4923/n76 ), .C(\DP_OP_665J1_134_4923/n77 ), .Y(
        \DP_OP_665J1_134_4923/n213 ) );
  NAND2XL \DP_OP_665J1_134_4923/U92  ( .A(N1447), .B(si_sel), .Y(
        \DP_OP_665J1_134_4923/n72 ) );
  NAND2XL \DP_OP_665J1_134_4923/U179  ( .A(N464), .B(\DP_OP_665J1_134_4923/I3 ), .Y(\DP_OP_665J1_134_4923/n140 ) );
  AOI22XL \DP_OP_665J1_134_4923/U181  ( .A0(n106), .A1(\C163/Z_1 ), .B0(
        \DP_OP_665J1_134_4923/I4 ), .B1(N580), .Y(\DP_OP_665J1_134_4923/n142 )
         );
  NAND3XL \DP_OP_665J1_134_4923/U178  ( .A(\DP_OP_665J1_134_4923/n141 ), .B(
        \DP_OP_665J1_134_4923/n140 ), .C(\DP_OP_665J1_134_4923/n142 ), .Y(
        \DP_OP_665J1_134_4923/n234 ) );
  NAND2XL \DP_OP_665J1_134_4923/U93  ( .A(\DP_OP_665J1_134_4923/n234 ), .B(
        \DP_OP_665J1_134_4923/I7 ), .Y(\DP_OP_665J1_134_4923/n73 ) );
  NAND2XL \DP_OP_665J1_134_4923/U94  ( .A(\DP_OP_665J1_134_4923/I10 ), .B(
        \U3/RSOP_657/C2/Z_1 ), .Y(\DP_OP_665J1_134_4923/n74 ) );
  NAND3XL \DP_OP_665J1_134_4923/U91  ( .A(\DP_OP_665J1_134_4923/n72 ), .B(
        \DP_OP_665J1_134_4923/n73 ), .C(\DP_OP_665J1_134_4923/n74 ), .Y(
        \DP_OP_665J1_134_4923/n214 ) );
  XOR2XL \DP_OP_665J1_134_4923/U2  ( .A(\DP_OP_665J1_134_4923/n232 ), .B(
        \C1/Z_19 ), .Y(\DP_OP_665J1_134_4923/n1 ) );
  XOR2XL \DP_OP_665J1_134_4923/U1  ( .A(\DP_OP_665J1_134_4923/n2 ), .B(
        \DP_OP_665J1_134_4923/n1 ), .Y(\C162/DATA3_19 ) );
  AND2XL \DP_OP_251J1_126_494/U12  ( .A(\C1/Z_0 ), .B(\DP_OP_251J1_126_494/I3 ), .Y(\DP_OP_251J1_126_494/n16 ) );
  AND2XL \DP_OP_251J1_126_494/U7  ( .A(\DP_OP_251J1_126_494/n27 ), .B(
        \DP_OP_251J1_126_494/I3 ), .Y(\DP_OP_251J1_126_494/n21 ) );
  DFFRX2 \write_cntr_reg/q_reg[10]  ( .D(n526), .CK(clk), .RN(n275), .Q(
        write_cntr[10]), .QN(n107) );
  DFFRX2 \work_cntr_reg[4]  ( .D(next_work_cntr[4]), .CK(clk), .RN(n274), .Q(
        work_cntr[4]), .QN(n180) );
  DFFRX4 \write_addr_reg/q_reg[16]  ( .D(n474), .CK(clk), .RN(n274), .Q(
        write_addr[16]), .QN(n248) );
  ADDHX1 \DP_OP_665J1_134_4923/U221  ( .A(write_addr[16]), .B(
        \DP_OP_665J1_134_4923/n178 ), .CO(\DP_OP_665J1_134_4923/n177 ), .S(
        N477) );
  ADDHX1 \DP_OP_665J1_134_4923/U209  ( .A(write_addr[16]), .B(
        \DP_OP_665J1_134_4923/n168 ), .CO(\DP_OP_665J1_134_4923/n167 ), .S(
        N593) );
  DFFRX2 \work_cntr_reg[10]  ( .D(next_work_cntr[10]), .CK(clk), .RN(n274), 
        .Q(work_cntr[10]), .QN(n183) );
  DFFRX2 \work_cntr_reg[19]  ( .D(next_work_cntr[19]), .CK(clk), .RN(n275), 
        .Q(work_cntr[19]), .QN(n212) );
  DFFRX2 \write_addr_reg/q_reg[14]  ( .D(n476), .CK(clk), .RN(n274), .Q(
        write_addr[14]), .QN(n246) );
  ADDHX1 \DP_OP_665J1_134_4923/U223  ( .A(write_addr[14]), .B(
        \DP_OP_665J1_134_4923/n180 ), .CO(\DP_OP_665J1_134_4923/n179 ), .S(
        N475) );
  ADDHX1 \DP_OP_665J1_134_4923/U211  ( .A(write_addr[14]), .B(
        \DP_OP_665J1_134_4923/n170 ), .CO(\DP_OP_665J1_134_4923/n169 ), .S(
        N591) );
  DFFRX2 \write_cntr_reg/q_reg[12]  ( .D(n524), .CK(clk), .RN(n709), .Q(
        write_cntr[12]), .QN(n211) );
  DFFRX2 \write_addr_reg/q_reg[11]  ( .D(n479), .CK(clk), .RN(n274), .Q(
        write_addr[11]), .QN(n245) );
  ADDHX1 \DP_OP_665J1_134_4923/U226  ( .A(write_addr[11]), .B(
        \DP_OP_665J1_134_4923/n183 ), .CO(\DP_OP_665J1_134_4923/n182 ), .S(
        N472) );
  ADDHX1 \DP_OP_665J1_134_4923/U214  ( .A(write_addr[11]), .B(
        \DP_OP_665J1_134_4923/n173 ), .CO(\DP_OP_665J1_134_4923/n172 ), .S(
        N588) );
  DFFRX2 \work_cntr_reg[12]  ( .D(next_work_cntr[12]), .CK(clk), .RN(n275), 
        .Q(work_cntr[12]), .QN(n215) );
  DFFRX2 \work_cntr_reg[9]  ( .D(next_work_cntr[9]), .CK(clk), .RN(n275), .Q(
        work_cntr[9]), .QN(n214) );
  DFFRX2 \work_cntr_reg[15]  ( .D(next_work_cntr[15]), .CK(clk), .RN(n275), 
        .Q(work_cntr[15]), .QN(n181) );
  DFFRX2 \work_cntr_reg[7]  ( .D(next_work_cntr[7]), .CK(clk), .RN(n274), .Q(
        work_cntr[7]), .QN(n176) );
  DFFRX4 \work_cntr_reg[14]  ( .D(next_work_cntr[14]), .CK(clk), .RN(n275), 
        .Q(work_cntr[14]), .QN(n219) );
  ADDHX1 \DP_OP_665J1_134_4923/U250  ( .A(N584), .B(
        \DP_OP_665J1_134_4923/n187 ), .CO(\DP_OP_665J1_134_4923/n203 ), .S(
        N468) );
  ADDHX1 \DP_OP_665J1_134_4923/U249  ( .A(N585), .B(
        \DP_OP_665J1_134_4923/n203 ), .CO(\DP_OP_665J1_134_4923/n202 ), .S(
        N469) );
  DFFRX2 \work_cntr_reg[0]  ( .D(next_work_cntr[0]), .CK(clk), .RN(n274), .Q(
        N85), .QN(n234) );
  DFFRX2 \write_addr_reg/q_reg[18]  ( .D(n472), .CK(clk), .RN(n274), .Q(
        write_addr[18]), .QN(n252) );
  DFFRX2 \work_cntr_reg[5]  ( .D(next_work_cntr[5]), .CK(clk), .RN(n274), .Q(
        work_cntr[5]), .QN(n168) );
  DFFRX2 \write_cntr_reg/q_reg[9]  ( .D(n527), .CK(clk), .RN(n274), .Q(
        write_cntr[9]), .QN(n203) );
  DFFRX2 \write_cntr_reg/q_reg[8]  ( .D(n534), .CK(clk), .RN(n274), .Q(
        write_cntr[8]), .QN(n173) );
  DFFRX4 \work_cntr_reg[2]  ( .D(next_work_cntr[2]), .CK(clk), .RN(n274), .Q(
        N2062), .QN(n167) );
  DFFRX4 \work_cntr_reg[3]  ( .D(next_work_cntr[3]), .CK(clk), .RN(n274), .Q(
        N2063), .QN(n179) );
  DFFRX2 \global_cntr_reg[9]  ( .D(n701), .CK(clk), .RN(n274), .Q(
        global_cntr[9]) );
  DFFRX2 \global_cntr_reg[2]  ( .D(next_glb_cntr[2]), .CK(clk), .RN(n709), .Q(
        global_cntr[2]), .QN(n161) );
  DFFRX4 \work_cntr_reg[8]  ( .D(next_work_cntr[8]), .CK(clk), .RN(n275), .Q(
        work_cntr[8]), .QN(n226) );
  DFFRX2 \work_cntr_reg[1]  ( .D(next_work_cntr[1]), .CK(clk), .RN(n274), .Q(
        N2061), .QN(n187) );
  DFFRX2 \write_addr_reg/q_reg[1]  ( .D(n489), .CK(clk), .RN(n709), .Q(N579), 
        .QN(n238) );
  DFFRX2 \write_addr_reg/q_reg[5]  ( .D(n485), .CK(clk), .RN(n274), .Q(N583), 
        .QN(n2310) );
  DFFRX2 \write_addr_reg/q_reg[13]  ( .D(n477), .CK(clk), .RN(n274), .Q(
        write_addr[13]), .QN(n166) );
  ADDHX1 \DP_OP_665J1_134_4923/U212  ( .A(write_addr[13]), .B(
        \DP_OP_665J1_134_4923/n171 ), .CO(\DP_OP_665J1_134_4923/n170 ), .S(
        N590) );
  ADDHX1 \DP_OP_665J1_134_4923/U224  ( .A(write_addr[13]), .B(
        \DP_OP_665J1_134_4923/n181 ), .CO(\DP_OP_665J1_134_4923/n180 ), .S(
        N474) );
  DFFRX2 \work_cntr_reg[16]  ( .D(next_work_cntr[16]), .CK(clk), .RN(n275), 
        .Q(work_cntr[16]), .QN(n182) );
  DFFRX2 \write_addr_reg/q_reg[9]  ( .D(n481), .CK(clk), .RN(n275), .Q(
        write_addr[9]), .QN(n244) );
  ADDHX1 \DP_OP_665J1_134_4923/U228  ( .A(write_addr[9]), .B(
        \DP_OP_665J1_134_4923/n202 ), .CO(\DP_OP_665J1_134_4923/n184 ), .S(
        N470) );
  DFFRX2 \write_addr_reg/q_reg[6]  ( .D(n484), .CK(clk), .RN(n709), .Q(N584), 
        .QN(n163) );
  DFFRX2 \work_cntr_reg[11]  ( .D(next_work_cntr[11]), .CK(clk), .RN(n275), 
        .Q(work_cntr[11]), .QN(n222) );
  DFFRX2 \write_addr_reg/q_reg[10]  ( .D(n480), .CK(clk), .RN(n274), .Q(
        write_addr[10]), .QN(n243) );
  ADDHX1 \DP_OP_665J1_134_4923/U227  ( .A(write_addr[10]), .B(
        \DP_OP_665J1_134_4923/n184 ), .CO(\DP_OP_665J1_134_4923/n183 ), .S(
        N471) );
  ADDHX1 \DP_OP_665J1_134_4923/U215  ( .A(write_addr[10]), .B(write_addr[9]), 
        .CO(\DP_OP_665J1_134_4923/n173 ), .S(N587) );
  DFFRX2 \write_addr_reg/q_reg[15]  ( .D(n475), .CK(clk), .RN(n274), .Q(
        write_addr[15]), .QN(n247) );
  ADDHX1 \DP_OP_665J1_134_4923/U222  ( .A(write_addr[15]), .B(
        \DP_OP_665J1_134_4923/n179 ), .CO(\DP_OP_665J1_134_4923/n178 ), .S(
        N476) );
  ADDHX1 \DP_OP_665J1_134_4923/U210  ( .A(write_addr[15]), .B(
        \DP_OP_665J1_134_4923/n169 ), .CO(\DP_OP_665J1_134_4923/n168 ), .S(
        N592) );
  DFFSX2 \state_reg[0]  ( .D(n14), .CK(clk), .SN(n275), .Q(n172), .QN(state[0]) );
  DFFRX2 \write_addr_reg/q_reg[2]  ( .D(n488), .CK(clk), .RN(n274), .Q(N580), 
        .QN(n235) );
  ADDHX1 \DP_OP_665J1_134_4923/U234  ( .A(N580), .B(N579), .CO(
        \DP_OP_665J1_134_4923/n190 ), .S(N464) );
  DFFRX2 \write_cntr_reg/q_reg[6]  ( .D(n529), .CK(clk), .RN(n709), .Q(
        write_cntr[6]), .QN(n209) );
  DFFRX2 \read_cntr_reg/q_reg[0]  ( .D(n519), .CK(clk), .RN(n274), .Q(
        read_cntr[0]), .QN(n170) );
  DFFRX2 \write_cntr_reg/q_reg[7]  ( .D(n528), .CK(clk), .RN(n709), .Q(
        write_cntr[7]), .QN(n1777) );
  DFFRX2 \work_cntr_reg[17]  ( .D(next_work_cntr[17]), .CK(clk), .RN(n275), 
        .Q(work_cntr[17]), .QN(n213) );
  DFFRX2 \write_addr_reg/q_reg[8]  ( .D(n482), .CK(clk), .RN(n275), .Q(
        write_addr[8]), .QN(n165) );
  DFFRX2 \work_cntr_reg[18]  ( .D(next_work_cntr[18]), .CK(clk), .RN(n275), 
        .Q(work_cntr[18]), .QN(n177) );
  DFFRX2 \write_addr_reg/q_reg[3]  ( .D(n487), .CK(clk), .RN(n274), .Q(N581), 
        .QN(n162) );
  ADDHX1 \DP_OP_665J1_134_4923/U253  ( .A(N581), .B(
        \DP_OP_665J1_134_4923/n190 ), .CO(\DP_OP_665J1_134_4923/n206 ), .S(
        N465) );
  ADDHX1 \DP_OP_665J1_134_4923/U252  ( .A(n272), .B(
        \DP_OP_665J1_134_4923/n206 ), .CO(\DP_OP_665J1_134_4923/n205 ), .S(
        N466) );
  ADDHX1 \DP_OP_665J1_134_4923/U231  ( .A(N583), .B(
        \DP_OP_665J1_134_4923/n205 ), .CO(\DP_OP_665J1_134_4923/n187 ), .S(
        N467) );
  DFFRX2 \write_addr_reg/q_reg[19]  ( .D(n471), .CK(clk), .RN(n274), .Q(
        write_addr[19]), .QN(n232) );
  DFFRX2 \write_cntr_reg/q_reg[11]  ( .D(n525), .CK(clk), .RN(n275), .Q(
        write_cntr[11]), .QN(n227) );
  DFFRX2 \work_cntr_reg[6]  ( .D(next_work_cntr[6]), .CK(clk), .RN(n274), .Q(
        work_cntr[6]), .QN(n178) );
  DFFRX2 \write_addr_reg/q_reg[7]  ( .D(n483), .CK(clk), .RN(n275), .Q(N585), 
        .QN(n241) );
  ADDHX1 \DP_OP_665J1_134_4923/U225  ( .A(write_addr[12]), .B(
        \DP_OP_665J1_134_4923/n182 ), .CO(\DP_OP_665J1_134_4923/n181 ), .S(
        N473) );
  ADDHX1 \DP_OP_665J1_134_4923/U213  ( .A(write_addr[12]), .B(
        \DP_OP_665J1_134_4923/n172 ), .CO(\DP_OP_665J1_134_4923/n171 ), .S(
        N589) );
  DFFRX4 \work_cntr_reg[13]  ( .D(next_work_cntr[13]), .CK(clk), .RN(n275), 
        .Q(work_cntr[13]), .QN(n221) );
  DFFRX2 \write_cntr_reg/q_reg[4]  ( .D(n535), .CK(clk), .RN(n275), .Q(
        write_cntr[4]) );
  ADDHX1 \DP_OP_665J1_134_4923/U220  ( .A(n271), .B(
        \DP_OP_665J1_134_4923/n177 ), .CO(\DP_OP_665J1_134_4923/n176 ), .S(
        N478) );
  ADDHX1 \DP_OP_665J1_134_4923/U219  ( .A(write_addr[18]), .B(
        \DP_OP_665J1_134_4923/n176 ), .CO(\DP_OP_665J1_134_4923/n175 ), .S(
        N479) );
  ADDHX1 \DP_OP_665J1_134_4923/U205  ( .A(fb_addr[0]), .B(
        \next_write_addr_w[0] ), .CO(\DP_OP_665J1_134_4923/n164 ), .S(N1446)
         );
  ADDHX1 \DP_OP_665J1_134_4923/U208  ( .A(n271), .B(
        \DP_OP_665J1_134_4923/n167 ), .CO(\DP_OP_665J1_134_4923/n166 ), .S(
        N594) );
  ADDHX1 \DP_OP_665J1_134_4923/U207  ( .A(write_addr[18]), .B(
        \DP_OP_665J1_134_4923/n166 ), .CO(\DP_OP_665J1_134_4923/n165 ), .S(
        N595) );
  ADDHX1 \DP_OP_665J1_134_4923/U206  ( .A(write_addr[19]), .B(
        \DP_OP_665J1_134_4923/n165 ), .CO(N597), .S(N596) );
  DFFRX2 \cr_read_cntr_reg/q_reg[6]  ( .D(n493), .CK(clk), .RN(n274), .Q(
        cr_read_cntr[6]) );
  DFFRX1 \state_reg[1]  ( .D(next_state[1]), .CK(clk), .RN(n709), .QN(n28) );
  DFFRX1 \global_cntr_reg[5]  ( .D(n705), .CK(clk), .RN(n709), .Q(
        global_cntr[5]), .QN(n630) );
  DFFRX1 \cr_read_cntr_reg/q_reg[0]  ( .D(n499), .CK(clk), .RN(n709), .Q(N1232), .QN(n4) );
  DFFRX1 \cr_read_cntr_reg/q_reg[3]  ( .D(n496), .CK(clk), .RN(n709), .Q(
        cr_read_cntr[3]) );
  DFFRX1 \global_cntr_reg[0]  ( .D(n236), .CK(clk), .RN(n709), .Q(
        global_cntr[0]), .QN(n236) );
  DFFRX1 \global_cntr_reg[1]  ( .D(next_glb_cntr[1]), .CK(clk), .RN(n709), .Q(
        global_cntr[1]), .QN(n204) );
  DFFRX1 \global_cntr_reg[3]  ( .D(n707), .CK(clk), .RN(n709), .Q(
        global_cntr[3]), .QN(n242) );
  DFFRX1 \global_cntr_reg[4]  ( .D(n706), .CK(clk), .RN(n709), .Q(
        global_cntr[4]), .QN(n190) );
  DFFRX1 \global_cntr_reg[6]  ( .D(n704), .CK(clk), .RN(n709), .Q(
        global_cntr[6]), .QN(n196) );
  DFFRX1 \global_cntr_reg[7]  ( .D(n703), .CK(clk), .RN(n709), .Q(
        global_cntr[7]), .QN(n194) );
  DFFRX1 \global_cntr_reg[8]  ( .D(n702), .CK(clk), .RN(n709), .Q(
        global_cntr[8]), .QN(n200) );
  DFFRX1 \global_cntr_reg[10]  ( .D(n700), .CK(clk), .RN(n709), .Q(
        global_cntr[10]), .QN(n197) );
  DFFRX1 \global_cntr_reg[11]  ( .D(n699), .CK(clk), .RN(n709), .Q(
        global_cntr[11]), .QN(n195) );
  DFFRX1 \global_cntr_reg[12]  ( .D(n698), .CK(clk), .RN(n709), .Q(
        global_cntr[12]), .QN(n198) );
  DFFRX1 \global_cntr_reg[13]  ( .D(n697), .CK(clk), .RN(n709), .Q(
        global_cntr[13]), .QN(n250) );
  DFFRX1 \global_cntr_reg[14]  ( .D(n696), .CK(clk), .RN(n709), .Q(
        global_cntr[14]), .QN(n201) );
  DFFRX1 \global_cntr_reg[15]  ( .D(n695), .CK(clk), .RN(n709), .Q(
        global_cntr[15]), .QN(n199) );
  DFFRX1 \global_cntr_reg[17]  ( .D(n693), .CK(clk), .RN(n709), .Q(
        global_cntr[17]), .QN(n202) );
  DFFRX1 \global_cntr_reg[16]  ( .D(n694), .CK(clk), .RN(n709), .Q(
        global_cntr[16]), .QN(n251) );
  DFFRX1 \global_cntr_reg[19]  ( .D(next_glb_cntr[19]), .CK(clk), .RN(n709), 
        .Q(global_cntr[19]), .QN(n255) );
  DFFRX1 \global_cntr_reg[18]  ( .D(n692), .CK(clk), .RN(n709), .Q(
        global_cntr[18]), .QN(n253) );
  DFFRX1 \state_reg[2]  ( .D(next_state[2]), .CK(clk), .RN(n709), .Q(state[2]), 
        .QN(n205) );
  DFFRX1 \curr_photo_reg[1]  ( .D(next_photo[1]), .CK(clk), .RN(n709), .Q(
        curr_photo[1]), .QN(n240) );
  DFFRX1 \curr_photo_reg[0]  ( .D(next_photo[0]), .CK(clk), .RN(n709), .Q(
        curr_photo[0]), .QN(n188) );
  DFFRX1 \read_cntr_reg/q_reg[1]  ( .D(n518), .CK(clk), .RN(n709), .Q(
        read_cntr[1]), .QN(n233) );
  DFFRX2 \write_addr_reg/q_reg[12]  ( .D(n478), .CK(clk), .RN(n709), .Q(
        write_addr[12]), .QN(n164) );
  ADDFX2 \DP_OP_251J1_126_494/U5  ( .A(\DP_OP_251J1_126_494/n5 ), .B(N32), 
        .CI(\DP_OP_251J1_126_494/n17 ), .CO(\DP_OP_251J1_126_494/n4 ), .S(
        N1236) );
  NOR2X1 U3 ( .A(n1674), .B(n1673), .Y(n1681) );
  CLKINVX1 U4 ( .A(next_cr_x[5]), .Y(n1223) );
  AOI2BB2X1 U5 ( .B0(n1272), .B1(n1271), .A0N(n1272), .A1N(n1268), .Y(n1276)
         );
  OR2X1 U6 ( .A(n375), .B(n934), .Y(n372) );
  CLKINVX1 U7 ( .A(n683), .Y(n1601) );
  MXI2X2 U8 ( .A(n401), .B(n402), .S0(n400), .Y(n421) );
  CLKINVX1 U9 ( .A(curr_photo_size[0]), .Y(n716) );
  NOR2X1 U10 ( .A(n202), .B(n296), .Y(n297) );
  NAND2X1 U11 ( .A(n295), .B(global_cntr[16]), .Y(n296) );
  NOR2X1 U12 ( .A(n294), .B(n199), .Y(n295) );
  OR2X1 U13 ( .A(n293), .B(n201), .Y(n294) );
  OR2X1 U14 ( .A(n729), .B(n196), .Y(n283) );
  NOR2X1 U15 ( .A(n1602), .B(n161), .Y(n708) );
  NAND2X1 U16 ( .A(n281), .B(global_cntr[5]), .Y(n729) );
  NOR2X1 U17 ( .A(n280), .B(n190), .Y(n281) );
  NOR3X1 U18 ( .A(n172), .B(n2328), .C(n738), .Y(n746) );
  AO21X1 U19 ( .A0(n689), .A1(\intadd_4/SUM[1] ), .B0(n1), .Y(n610) );
  OAI21XL U20 ( .A0(n265), .A1(n243), .B0(n345), .Y(n1) );
  AND2X2 U21 ( .A(global_cntr[8]), .B(n284), .Y(n285) );
  OAI2BB2XL U22 ( .B0(n1326), .B1(n1324), .A0N(n1326), .A1N(n1324), .Y(n2) );
  OR2X1 U23 ( .A(n4), .B(n2334), .Y(n3) );
  OR2X1 U24 ( .A(n259), .B(n2334), .Y(n5) );
  OR2X1 U25 ( .A(n257), .B(n2334), .Y(n6) );
  OR2X1 U26 ( .A(n8), .B(n2334), .Y(n7) );
  XNOR2X1 U27 ( .A(\DP_OP_251J1_126_494/n1 ), .B(\DP_OP_251J1_126_494/n21 ), 
        .Y(n8) );
  AOI21X1 U28 ( .A0(n676), .A1(\C162/DATA3_3 ), .B0(n10), .Y(\im_a[3]_BAR ) );
  AO22X1 U29 ( .A0(n269), .A1(N1449), .B0(n268), .B1(global_cntr[3]), .Y(n10)
         );
  AOI21X1 U30 ( .A0(n676), .A1(\C162/DATA3_4 ), .B0(n12), .Y(\im_a[4]_BAR ) );
  AO22X1 U31 ( .A0(n269), .A1(N1450), .B0(n268), .B1(global_cntr[4]), .Y(n12)
         );
  AOI21X1 U32 ( .A0(n676), .A1(\C162/DATA3_5 ), .B0(n15), .Y(\im_a[5]_BAR ) );
  AO22X1 U33 ( .A0(n269), .A1(N1451), .B0(n268), .B1(global_cntr[5]), .Y(n15)
         );
  AOI21X1 U34 ( .A0(n676), .A1(\C162/DATA3_6 ), .B0(n17), .Y(\im_a[6]_BAR ) );
  AO22X1 U35 ( .A0(n269), .A1(N1452), .B0(n268), .B1(global_cntr[6]), .Y(n17)
         );
  AOI21X1 U36 ( .A0(n676), .A1(\C162/DATA3_7 ), .B0(n19), .Y(\im_a[7]_BAR ) );
  AO22X1 U37 ( .A0(n269), .A1(N1453), .B0(n268), .B1(global_cntr[7]), .Y(n19)
         );
  AOI21X1 U38 ( .A0(n676), .A1(\C162/DATA3_8 ), .B0(n21), .Y(\im_a[8]_BAR ) );
  AO22X1 U39 ( .A0(n269), .A1(N1454), .B0(n268), .B1(global_cntr[8]), .Y(n21)
         );
  AOI21X1 U40 ( .A0(n676), .A1(\C162/DATA3_9 ), .B0(n23), .Y(\im_a[9]_BAR ) );
  AO22X1 U41 ( .A0(n269), .A1(N1455), .B0(n268), .B1(global_cntr[9]), .Y(n23)
         );
  AOI21X1 U42 ( .A0(n676), .A1(\C162/DATA3_10 ), .B0(n25), .Y(\im_a[10]_BAR )
         );
  AO22X1 U43 ( .A0(n269), .A1(N1456), .B0(n268), .B1(global_cntr[10]), .Y(n25)
         );
  AOI21X1 U44 ( .A0(n676), .A1(\C162/DATA3_11 ), .B0(n27), .Y(\im_a[11]_BAR )
         );
  AO22X1 U45 ( .A0(n269), .A1(N1457), .B0(n268), .B1(global_cntr[11]), .Y(n27)
         );
  AOI21X1 U46 ( .A0(n676), .A1(\C162/DATA3_12 ), .B0(n30), .Y(\im_a[12]_BAR )
         );
  AO22X1 U47 ( .A0(n269), .A1(N1458), .B0(n268), .B1(global_cntr[12]), .Y(n30)
         );
  AOI21X1 U48 ( .A0(n676), .A1(\C162/DATA3_13 ), .B0(n32), .Y(\im_a[13]_BAR )
         );
  AO22X1 U49 ( .A0(n269), .A1(N1459), .B0(n268), .B1(global_cntr[13]), .Y(n32)
         );
  AOI21X1 U50 ( .A0(n676), .A1(\C162/DATA3_14 ), .B0(n34), .Y(\im_a[14]_BAR )
         );
  AO22X1 U51 ( .A0(n269), .A1(N1460), .B0(n268), .B1(global_cntr[14]), .Y(n34)
         );
  AOI21X1 U52 ( .A0(n676), .A1(\C162/DATA3_15 ), .B0(n36), .Y(\im_a[15]_BAR )
         );
  AO22X1 U53 ( .A0(n269), .A1(N1461), .B0(n268), .B1(global_cntr[15]), .Y(n36)
         );
  AOI21X1 U54 ( .A0(n676), .A1(\C162/DATA3_16 ), .B0(n38), .Y(\im_a[16]_BAR )
         );
  AO22X1 U55 ( .A0(n269), .A1(N1462), .B0(n268), .B1(global_cntr[16]), .Y(n38)
         );
  AOI21X1 U56 ( .A0(n676), .A1(\C162/DATA3_18 ), .B0(n40), .Y(\im_a[18]_BAR )
         );
  AO22X1 U57 ( .A0(n269), .A1(N1464), .B0(n268), .B1(global_cntr[18]), .Y(n40)
         );
  OR2X2 U58 ( .A(state[2]), .B(n28), .Y(n2328) );
  NAND2X1 U59 ( .A(global_cntr[2]), .B(n1602), .Y(n1516) );
  NAND2X1 U60 ( .A(state[2]), .B(n28), .Y(n742) );
  CLKINVX1 U61 ( .A(n2120), .Y(n1922) );
  NOR2X1 U62 ( .A(n1353), .B(n1761), .Y(n2289) );
  AOI2BB1X1 U63 ( .A0N(write_cntr[12]), .A1N(n1521), .B0(n230), .Y(n1532) );
  OAI2BB1X1 U64 ( .A0N(n384), .A1N(\s_1[3] ), .B0(n941), .Y(n392) );
  NAND2BX1 U65 ( .AN(n313), .B(n926), .Y(n406) );
  OAI2BB1X1 U66 ( .A0N(n302), .A1N(h_1[3]), .B0(n919), .Y(n311) );
  NAND2BX1 U67 ( .AN(n403), .B(n458), .Y(n450) );
  OAI22XL U68 ( .A0(n1304), .A1(n1355), .B0(n164), .B1(n265), .Y(n41) );
  AOI211X1 U69 ( .A0(\intadd_4/SUM[3] ), .A1(n689), .B0(n1305), .C0(n41), .Y(
        n42) );
  CLKINVX1 U70 ( .A(n42), .Y(n595) );
  NAND2BX1 U71 ( .AN(n1522), .B(write_cntr[14]), .Y(n1531) );
  CLKINVX1 U72 ( .A(\m_1[3] ), .Y(n43) );
  NAND2X1 U73 ( .A(n415), .B(n411), .Y(n44) );
  AOI211X1 U74 ( .A0(n382), .A1(n44), .B0(n412), .C0(n465), .Y(n45) );
  CLKINVX1 U75 ( .A(\s_1[3] ), .Y(n46) );
  AO22X1 U76 ( .A0(n420), .A1(n421), .B0(n419), .B1(n418), .Y(n47) );
  OAI22XL U77 ( .A0(n450), .A1(n46), .B0(n440), .B1(n47), .Y(n48) );
  AOI211X1 U78 ( .A0(n463), .A1(h_1[3]), .B0(n45), .C0(n48), .Y(n49) );
  OA21XL U79 ( .A0(n926), .A1(n410), .B0(n409), .Y(n50) );
  NAND2X1 U80 ( .A(n454), .B(n430), .Y(n51) );
  NAND2X1 U81 ( .A(n50), .B(n51), .Y(n52) );
  OAI211X1 U82 ( .A0(n50), .A1(n51), .B0(n464), .C0(n52), .Y(n53) );
  OAI211X1 U83 ( .A0(n466), .A1(n43), .B0(n49), .C0(n53), .Y(\C1/Z_3 ) );
  AO22X1 U84 ( .A0(N474), .A1(\DP_OP_665J1_134_4923/I2 ), .B0(
        \DP_OP_665J1_134_4923/I3 ), .B1(\DP_OP_665J1_134_4923/n263 ), .Y(n54)
         );
  AOI22X1 U85 ( .A0(N590), .A1(n267), .B0(N474), .B1(n567), .Y(n55) );
  NAND2X1 U86 ( .A(write_addr[13]), .B(n568), .Y(n56) );
  OAI211X1 U87 ( .A0(n571), .A1(n596), .B0(n55), .C0(n56), .Y(n57) );
  AO22X1 U88 ( .A0(\DP_OP_665J1_134_4923/I4 ), .A1(N590), .B0(n106), .B1(n57), 
        .Y(n58) );
  OAI21XL U89 ( .A0(n54), .A1(n58), .B0(\DP_OP_665J1_134_4923/I7 ), .Y(
        \DP_OP_665J1_134_4923/n43 ) );
  AO21X1 U90 ( .A0(n244), .A1(n1295), .B0(n1294), .Y(n59) );
  AO21X1 U91 ( .A0(n1297), .A1(n59), .B0(n1327), .Y(n60) );
  OAI222XL U92 ( .A0(n60), .A1(n1296), .B0(n59), .B1(n1355), .C0(n265), .C1(
        n244), .Y(n61) );
  AOI2BB1X1 U93 ( .A0N(n1353), .A1N(\intadd_3/SUM[6] ), .B0(n61), .Y(n612) );
  OAI2BB1X1 U94 ( .A0N(n1533), .A1N(n1532), .B0(n1531), .Y(n1580) );
  OAI2BB1X1 U95 ( .A0N(n392), .A1N(n393), .B0(n394), .Y(n395) );
  AO21X1 U96 ( .A0(n62), .A1(h_1[1]), .B0(n925), .Y(n409) );
  CLKINVX1 U97 ( .A(curr_time[18]), .Y(n62) );
  AO22X1 U98 ( .A0(N477), .A1(\DP_OP_665J1_134_4923/I2 ), .B0(
        \DP_OP_665J1_134_4923/I3 ), .B1(\DP_OP_665J1_134_4923/n266 ), .Y(n63)
         );
  AOI22X1 U99 ( .A0(N593), .A1(n267), .B0(N477), .B1(n567), .Y(n64) );
  NAND2X1 U100 ( .A(write_addr[16]), .B(n568), .Y(n65) );
  OAI211X1 U101 ( .A0(n571), .A1(n586), .B0(n64), .C0(n65), .Y(n66) );
  AO22X1 U102 ( .A0(\DP_OP_665J1_134_4923/I4 ), .A1(N593), .B0(n106), .B1(n66), 
        .Y(n67) );
  OAI21XL U103 ( .A0(n63), .A1(n67), .B0(\DP_OP_665J1_134_4923/I7 ), .Y(
        \DP_OP_665J1_134_4923/n34 ) );
  AO21X1 U104 ( .A0(\DP_OP_251J1_126_494/n24 ), .A1(\DP_OP_251J1_126_494/I3 ), 
        .B0(\DP_OP_251J1_126_494/I2 ), .Y(n68) );
  AND2X1 U105 ( .A(\DP_OP_251J1_126_494/n4 ), .B(n68), .Y(
        \DP_OP_251J1_126_494/n3 ) );
  AOI2BB2X1 U106 ( .B0(\DP_OP_251J1_126_494/n4 ), .B1(n68), .A0N(
        \DP_OP_251J1_126_494/n4 ), .A1N(n68), .Y(N1237) );
  CLKINVX1 U107 ( .A(n702), .Y(n69) );
  OAI21XL U108 ( .A0(n734), .A1(n69), .B0(n730), .Y(n70) );
  NAND3XL U109 ( .A(global_cntr[11]), .B(n700), .C(n70), .Y(n71) );
  CLKINVX1 U110 ( .A(n694), .Y(n72) );
  AOI211X1 U111 ( .A0(n735), .A1(n71), .B0(n202), .C0(n72), .Y(n73) );
  OR3X1 U112 ( .A(n692), .B(next_glb_cntr[19]), .C(n73), .Y(n738) );
  CLKINVX1 U113 ( .A(n1328), .Y(n74) );
  AOI2BB2X1 U114 ( .B0(n1329), .B1(n1328), .A0N(n1329), .A1N(n271), .Y(n75) );
  OAI222XL U115 ( .A0(n74), .A1(n1355), .B0(n75), .B1(n1327), .C0(n231), .C1(
        n265), .Y(n76) );
  CLKINVX1 U116 ( .A(n76), .Y(n582) );
  NOR2X1 U117 ( .A(n1002), .B(n1264), .Y(n77) );
  XNOR2X1 U118 ( .A(n77), .B(n828), .Y(n844) );
  NAND2X1 U119 ( .A(n768), .B(next_cr_x[6]), .Y(n78) );
  XNOR2X1 U120 ( .A(n78), .B(n769), .Y(n967) );
  OAI2BB1X1 U121 ( .A0N(n1546), .A1N(n1547), .B0(n1545), .Y(n1579) );
  OAI2BB1X1 U122 ( .A0N(n316), .A1N(\m_1[3] ), .B0(n931), .Y(n374) );
  CLKINVX1 U123 ( .A(curr_time[4]), .Y(n79) );
  NAND2X1 U124 ( .A(n387), .B(n392), .Y(n80) );
  OAI211X1 U125 ( .A0(n941), .A1(n79), .B0(n942), .C0(n80), .Y(n394) );
  CLKINVX1 U126 ( .A(curr_time[20]), .Y(n81) );
  NAND2X1 U127 ( .A(n305), .B(n311), .Y(n82) );
  OAI211X1 U128 ( .A0(n919), .A1(n81), .B0(n922), .C0(n82), .Y(n310) );
  AO22X1 U129 ( .A0(N481), .A1(\DP_OP_665J1_134_4923/I2 ), .B0(
        \DP_OP_665J1_134_4923/I3 ), .B1(\DP_OP_665J1_134_4923/n270 ), .Y(n83)
         );
  AO22X1 U130 ( .A0(N597), .A1(n267), .B0(N481), .B1(n567), .Y(n84) );
  AO22X1 U131 ( .A0(\DP_OP_665J1_134_4923/I4 ), .A1(N597), .B0(n106), .B1(n84), 
        .Y(n85) );
  OAI21XL U132 ( .A0(n83), .A1(n85), .B0(\DP_OP_665J1_134_4923/I7 ), .Y(
        \DP_OP_665J1_134_4923/n22 ) );
  AO21X1 U133 ( .A0(\DP_OP_251J1_126_494/n25 ), .A1(\DP_OP_251J1_126_494/I3 ), 
        .B0(\DP_OP_251J1_126_494/I2 ), .Y(n86) );
  AND2X1 U134 ( .A(\DP_OP_251J1_126_494/n3 ), .B(n86), .Y(
        \DP_OP_251J1_126_494/n2 ) );
  AOI2BB2X1 U135 ( .B0(\DP_OP_251J1_126_494/n3 ), .B1(n86), .A0N(
        \DP_OP_251J1_126_494/n3 ), .A1N(n86), .Y(N1238) );
  AO21X1 U136 ( .A0(n2340), .A1(n2291), .B0(n2290), .Y(n365) );
  AOI32X1 U137 ( .A0(n1615), .A1(n1617), .A2(n1620), .B0(n1619), .B1(n1617), 
        .Y(n1631) );
  OAI2BB1X1 U138 ( .A0N(n126), .A1N(n848), .B0(n842), .Y(n1269) );
  CLKINVX1 U139 ( .A(curr_time[12]), .Y(n87) );
  NAND2X1 U140 ( .A(n319), .B(n374), .Y(n88) );
  OAI211X1 U141 ( .A0(n931), .A1(n87), .B0(n934), .C0(n88), .Y(n373) );
  OAI2BB1X1 U142 ( .A0N(n1561), .A1N(n1560), .B0(n1559), .Y(n1578) );
  AOI2BB1X1 U143 ( .A0N(n1688), .A1N(n1697), .B0(n1681), .Y(n89) );
  NAND2X1 U144 ( .A(n1678), .B(n1675), .Y(n90) );
  AOI2BB2X1 U145 ( .B0(n89), .B1(n90), .A0N(n89), .A1N(n90), .Y(n1685) );
  OAI2BB1X1 U146 ( .A0N(n399), .A1N(n400), .B0(n395), .Y(n438) );
  CLKINVX1 U147 ( .A(n711), .Y(n91) );
  AOI2BB2X1 U148 ( .B0(n91), .B1(n927), .A0N(n91), .A1N(h_1[1]), .Y(n928) );
  OR2X1 U149 ( .A(write_addr[9]), .B(\DP_OP_665J1_134_4923/n202 ), .Y(n92) );
  AOI2BB2X1 U150 ( .B0(write_addr[10]), .B1(n92), .A0N(write_addr[10]), .A1N(
        n92), .Y(\DP_OP_665J1_134_4923/n260 ) );
  AND2X1 U151 ( .A(write_addr[10]), .B(n92), .Y(\DP_OP_665J1_134_4923/n200 )
         );
  NAND2X1 U152 ( .A(\next_cr_y[0] ), .B(next_cr_x[5]), .Y(n93) );
  AOI2BB2X1 U153 ( .B0(next_cr_x[6]), .B1(n93), .A0N(next_cr_x[6]), .A1N(n93), 
        .Y(n94) );
  AOI2BB2X1 U154 ( .B0(n1240), .B1(n94), .A0N(n1240), .A1N(n94), .Y(
        \intadd_4/SUM[0] ) );
  CLKINVX1 U155 ( .A(next_cr_x[6]), .Y(n95) );
  AOI222XL U156 ( .A0(n1240), .A1(n93), .B0(n1240), .B1(n95), .C0(n93), .C1(
        n95), .Y(\intadd_4/n4 ) );
  NOR2X1 U157 ( .A(n594), .B(n641), .Y(n96) );
  OAI22XL U158 ( .A0(n246), .A1(n648), .B0(n164), .B1(n649), .Y(n97) );
  AOI211X1 U159 ( .A0(n595), .A1(n645), .B0(n96), .C0(n97), .Y(n98) );
  OAI22XL U160 ( .A0(n276), .A1(n201), .B0(n660), .B1(n98), .Y(n99) );
  NAND2X1 U161 ( .A(\DP_OP_665J1_134_4923/I10 ), .B(n99), .Y(
        \DP_OP_665J1_134_4923/n35 ) );
  AOI2BB2X1 U162 ( .B0(write_addr[19]), .B1(fb_addr[19]), .A0N(write_addr[19]), 
        .A1N(fb_addr[19]), .Y(n100) );
  AOI2BB2X1 U163 ( .B0(\DP_OP_665J1_134_4923/n146 ), .B1(n100), .A0N(
        \DP_OP_665J1_134_4923/n146 ), .A1N(n100), .Y(N1465) );
  AO21X1 U164 ( .A0(\DP_OP_251J1_126_494/n26 ), .A1(\DP_OP_251J1_126_494/I3 ), 
        .B0(\DP_OP_251J1_126_494/I2 ), .Y(n101) );
  AND2X1 U165 ( .A(\DP_OP_251J1_126_494/n2 ), .B(n101), .Y(
        \DP_OP_251J1_126_494/n1 ) );
  AOI2BB2X1 U166 ( .B0(\DP_OP_251J1_126_494/n2 ), .B1(n101), .A0N(
        \DP_OP_251J1_126_494/n2 ), .A1N(n101), .Y(N1239) );
  CLKINVX1 U167 ( .A(write_cntr[12]), .Y(n102) );
  OAI31XL U168 ( .A0(n755), .A1(n270), .A2(n102), .B0(n230), .Y(n103) );
  OAI21XL U169 ( .A0(n753), .A1(n270), .B0(n885), .Y(n104) );
  NAND2X1 U170 ( .A(n103), .B(n104), .Y(n787) );
  OR2X1 U171 ( .A(n277), .B(n2284), .Y(n1308) );
  OAI21XL U172 ( .A0(n295), .A1(global_cntr[16]), .B0(n296), .Y(n105) );
  NOR2X1 U173 ( .A(n731), .B(n105), .Y(n694) );
  NOR2BX1 U174 ( .AN(n1602), .B(n279), .Y(next_glb_cntr[1]) );
  OAI2BB2XL U175 ( .B0(n686), .B1(n2307), .A0N(n273), .A1N(N580), .Y(n488) );
  INVXL U176 ( .A(n654), .Y(n124) );
  AOI211X1 U177 ( .A0(n1065), .A1(n1245), .B0(n1064), .C0(n1063), .Y(n654) );
  OR3X4 U178 ( .A(n685), .B(n684), .C(n572), .Y(n106) );
  OR2X1 U179 ( .A(\intadd_3/B[0] ), .B(n1054), .Y(n1208) );
  AO21X1 U180 ( .A0(n690), .A1(n1764), .B0(n2290), .Y(n773) );
  OAI211X1 U181 ( .A0(n1074), .A1(n1073), .B0(n1072), .C0(n1071), .Y(n1079) );
  OA21X2 U182 ( .A0(n265), .A1(n247), .B0(n1321), .Y(n108) );
  NOR2X2 U183 ( .A(n277), .B(n1954), .Y(next_work_cntr[9]) );
  NOR2X2 U184 ( .A(n277), .B(n1958), .Y(next_work_cntr[15]) );
  NOR2X2 U185 ( .A(n277), .B(n1956), .Y(next_work_cntr[7]) );
  NOR2X2 U186 ( .A(n277), .B(n1951), .Y(next_work_cntr[14]) );
  INVX6 U187 ( .A(reset), .Y(n709) );
  BUFX4 U188 ( .A(n709), .Y(n275) );
  NAND2X2 U189 ( .A(n1212), .B(n1204), .Y(\next_cr_y[0] ) );
  OAI21X1 U190 ( .A0(n2286), .A1(n2285), .B0(n2284), .Y(n2291) );
  NOR2X1 U191 ( .A(n2223), .B(n2222), .Y(n2234) );
  OAI21X1 U192 ( .A0(n113), .A1(n860), .B0(n859), .Y(n867) );
  AND3X1 U193 ( .A(n266), .B(n332), .C(n1765), .Y(n2341) );
  NAND2X1 U194 ( .A(n2195), .B(n2210), .Y(n2219) );
  OAI22X1 U195 ( .A0(n1756), .A1(n1741), .B0(n1740), .B1(n1750), .Y(
        expand_sel[2]) );
  OAI21X1 U196 ( .A0(n1911), .A1(n1920), .B0(n1917), .Y(n1912) );
  OR2X4 U197 ( .A(n266), .B(n681), .Y(n660) );
  INVX1 U198 ( .A(n1184), .Y(n109) );
  OAI22X1 U199 ( .A0(n962), .A1(n995), .B0(n1779), .B1(n1230), .Y(n963) );
  OAI21X1 U200 ( .A0(n971), .A1(n970), .B0(n969), .Y(n1003) );
  INVXL U201 ( .A(n1825), .Y(n110) );
  AOI2BB2X2 U202 ( .B0(n1741), .B1(n1607), .A0N(n1609), .A1N(N85), .Y(
        expand_sel[0]) );
  NOR2BX1 U203 ( .AN(en_so), .B(n1764), .Y(n1765) );
  NAND2X1 U204 ( .A(curr_time[15]), .B(n930), .Y(n319) );
  NAND2X1 U205 ( .A(curr_time[7]), .B(n940), .Y(n387) );
  NAND2X2 U206 ( .A(global_cntr[1]), .B(global_cntr[0]), .Y(n1602) );
  OA21XL U207 ( .A0(n1211), .A1(n1218), .B0(n1210), .Y(n1337) );
  OA21XL U208 ( .A0(n1207), .A1(n1224), .B0(\intadd_3/CI ), .Y(n1338) );
  AOI32X1 U209 ( .A0(n2293), .A1(n682), .A2(cr_read_cntr[3]), .B0(n2299), .B1(
        n682), .Y(n2295) );
  OAI211X1 U210 ( .A0(n2257), .A1(n2256), .B0(n2263), .C0(n2255), .Y(n2261) );
  OAI31X1 U211 ( .A0(n2248), .A1(n2251), .A2(n2245), .B0(n2242), .Y(n2247) );
  NAND2X6 U212 ( .A(n2340), .B(im_wen_n), .Y(n2314) );
  OR2XL U213 ( .A(n858), .B(n857), .Y(n861) );
  OAI31X1 U214 ( .A0(n1751), .A1(n1750), .A2(n179), .B0(n1749), .Y(
        expand_sel[3]) );
  NAND2X4 U215 ( .A(n276), .B(n660), .Y(\DP_OP_665J1_134_4923/I10 ) );
  NAND3X6 U216 ( .A(n266), .B(n276), .C(n2334), .Y(n676) );
  OR2X1 U217 ( .A(n149), .B(n150), .Y(n148) );
  OA21XL U218 ( .A0(n1897), .A1(n1896), .B0(n1895), .Y(n1904) );
  OAI31X1 U219 ( .A0(n823), .A1(n994), .A2(n822), .B0(n821), .Y(n833) );
  OAI221X1 U220 ( .A0(work_cntr[5]), .A1(n2057), .B0(n1721), .B1(n2057), .C0(
        n1724), .Y(n1722) );
  OA21XL U221 ( .A0(n1483), .A1(n1482), .B0(n1481), .Y(n1491) );
  OA21XL U222 ( .A0(n1881), .A1(n1880), .B0(n1879), .Y(n1887) );
  OAI31X1 U223 ( .A0(n1251), .A1(n1254), .A2(n184), .B0(n1250), .Y(n1255) );
  OA21XL U224 ( .A0(n1914), .A1(n1180), .B0(n1185), .Y(n1184) );
  AOI222X1 U225 ( .A0(n2100), .A1(n2099), .B0(n2100), .B1(n2102), .C0(n2099), 
        .C1(n2098), .Y(n2101) );
  OAI211X1 U226 ( .A0(N2063), .A1(n2120), .B0(n1180), .C0(n1179), .Y(n1185) );
  OAI211X1 U227 ( .A0(n933), .A1(n466), .B0(n434), .C0(n433), .Y(\C1/Z_2 ) );
  OAI211X1 U228 ( .A0(n457), .A1(n466), .B0(n456), .C0(n455), .Y(\C1/Z_0 ) );
  OAI31X1 U229 ( .A0(n1457), .A1(work_cntr[6]), .A2(n1456), .B0(n1455), .Y(
        n1463) );
  NOR2X2 U230 ( .A(n791), .B(n795), .Y(n1248) );
  AOI211X1 U231 ( .A0(n1674), .A1(n1678), .B0(n1670), .C0(n1679), .Y(n1676) );
  AO22XL U232 ( .A0(n767), .A1(n783), .B0(n773), .B1(write_cntr[8]), .Y(n1772)
         );
  OA21XL U233 ( .A0(n1833), .A1(n1832), .B0(n1831), .Y(n1842) );
  NAND2BX2 U234 ( .AN(n277), .B(n299), .Y(n1353) );
  OA21XL U235 ( .A0(n1824), .A1(n1818), .B0(n1960), .Y(n1825) );
  OA21X4 U236 ( .A0(n205), .A1(next_state[2]), .B0(n744), .Y(n2340) );
  CLKINVX1 U237 ( .A(n14), .Y(n1059) );
  OAI31X1 U238 ( .A0(n298), .A1(n2328), .A2(n172), .B0(n737), .Y(next_state[2]) );
  OA21XL U239 ( .A0(n1411), .A1(n1410), .B0(n1409), .Y(n1415) );
  OAI31X1 U240 ( .A0(global_cntr[0]), .A1(n204), .A2(n161), .B0(n2279), .Y(
        n745) );
  OAI2BB1X4 U241 ( .A0N(read_cntr[1]), .A1N(n1365), .B0(n508), .Y(n567) );
  OR2X1 U242 ( .A(n152), .B(n153), .Y(n151) );
  NOR3XL U243 ( .A(n236), .B(n1516), .C(n1604), .Y(N2644) );
  NOR4X1 U244 ( .A(global_cntr[3]), .B(global_cntr[4]), .C(n1514), .D(n1513), 
        .Y(n1515) );
  BUFX8 U245 ( .A(n275), .Y(n274) );
  CLKINVX1 U246 ( .A(curr_photo_size[1]), .Y(n367) );
  INVX3 U247 ( .A(n961), .Y(n1779) );
  NAND2X1 U248 ( .A(n1581), .B(n1518), .Y(n1768) );
  NAND2X1 U249 ( .A(n1686), .B(n1685), .Y(n1699) );
  CLKINVX1 U250 ( .A(n1696), .Y(n1686) );
  NAND2X1 U251 ( .A(n181), .B(n1076), .Y(n1075) );
  CLKINVX1 U252 ( .A(n1077), .Y(n1076) );
  OAI21X1 U253 ( .A0(n1429), .A1(n1424), .B0(n183), .Y(n1430) );
  OAI21X1 U254 ( .A0(n1267), .A1(n1260), .B0(n1266), .Y(n1265) );
  OAI21X1 U255 ( .A0(n270), .A1(n782), .B0(n885), .Y(n781) );
  OAI21X1 U256 ( .A0(n232), .A1(n1055), .B0(n1056), .Y(n1058) );
  OAI21X1 U257 ( .A0(n2045), .A1(n2044), .B0(n2043), .Y(n2048) );
  OAI21X1 U258 ( .A0(n2080), .A1(n2079), .B0(n2078), .Y(n2083) );
  OAI21X1 U259 ( .A0(n2028), .A1(n2027), .B0(n2026), .Y(n2031) );
  CLKINVX1 U260 ( .A(n2021), .Y(n2028) );
  OAI21X1 U261 ( .A0(n1924), .A1(n1928), .B0(n1923), .Y(n1931) );
  OAI21X1 U262 ( .A0(n1155), .A1(n1154), .B0(n1153), .Y(n1162) );
  AOI211X1 U263 ( .A0(n2159), .A1(n2163), .B0(n2158), .C0(n2164), .Y(n2161) );
  NOR2X1 U264 ( .A(n2152), .B(n2151), .Y(n2158) );
  OAI22X1 U265 ( .A0(n2036), .A1(n2044), .B0(n2035), .B1(n2034), .Y(n2046) );
  OAI22X1 U266 ( .A0(n2072), .A1(n2079), .B0(n2071), .B1(n2070), .Y(n2081) );
  AOI2BB2X2 U267 ( .B0(write_cntr[10]), .B1(n1525), .A0N(write_cntr[10]), 
        .A1N(n1525), .Y(n1542) );
  OAI211X1 U268 ( .A0(n449), .A1(n466), .B0(n448), .C0(n447), .Y(\C1/Z_1 ) );
  NAND2X2 U269 ( .A(n460), .B(n1767), .Y(n466) );
  INVXL U270 ( .A(N480), .Y(n111) );
  INVXL U271 ( .A(n111), .Y(n112) );
  OAI22X1 U272 ( .A0(n960), .A1(n959), .B0(n968), .B1(n958), .Y(n1005) );
  NOR3X1 U273 ( .A(n212), .B(n177), .C(work_cntr[17]), .Y(n1375) );
  OAI31X1 U274 ( .A0(n1031), .A1(n1046), .A2(n1052), .B0(n1049), .Y(n1051) );
  NOR3BX1 U275 ( .AN(n1039), .B(n1042), .C(n1771), .Y(n1031) );
  NOR3BX1 U276 ( .AN(n2151), .B(n2155), .C(n2164), .Y(n2156) );
  AOI2BB2X2 U277 ( .B0(n2001), .B1(n2000), .A0N(n2001), .A1N(n1999), .Y(n2011)
         );
  BUFX4 U278 ( .A(n566), .Y(n267) );
  NOR2X2 U279 ( .A(n325), .B(n663), .Y(n664) );
  NOR2X1 U280 ( .A(n212), .B(n1781), .Y(n1784) );
  NAND2X1 U281 ( .A(n213), .B(n177), .Y(n1781) );
  CLKINVX1 U282 ( .A(n861), .Y(n113) );
  NOR2X1 U283 ( .A(n1999), .B(n1998), .Y(n2009) );
  NOR2X1 U284 ( .A(n213), .B(n1783), .Y(n956) );
  OAI21X1 U285 ( .A0(n1981), .A1(n182), .B0(n1982), .Y(n1619) );
  OAI21X1 U286 ( .A0(n1151), .A1(n1159), .B0(n1150), .Y(n1166) );
  OAI21X1 U287 ( .A0(curr_time[7]), .A1(n714), .B0(n939), .Y(n941) );
  CLKINVX1 U288 ( .A(n440), .Y(n462) );
  NAND2X1 U289 ( .A(n14), .B(n2278), .Y(n2284) );
  CLKINVX1 U290 ( .A(n2281), .Y(n2278) );
  OAI31X1 U291 ( .A0(n1401), .A1(work_cntr[13]), .A2(n1400), .B0(n1399), .Y(
        n1407) );
  NAND2X1 U292 ( .A(n1392), .B(n1393), .Y(n1401) );
  OAI31X1 U293 ( .A0(n1473), .A1(work_cntr[4]), .A2(n1472), .B0(n1471), .Y(
        n1479) );
  NAND2X1 U294 ( .A(n1464), .B(n1465), .Y(n1473) );
  OAI31X1 U295 ( .A0(n1852), .A1(n1851), .A2(n1850), .B0(n1849), .Y(n1856) );
  NAND2X1 U296 ( .A(n1843), .B(n1845), .Y(n1852) );
  OAI31X1 U297 ( .A0(n1886), .A1(n1885), .A2(n1884), .B0(n1883), .Y(n1892) );
  NAND2X1 U298 ( .A(n1875), .B(n1876), .Y(n1886) );
  OAI31X1 U299 ( .A0(n1868), .A1(n1867), .A2(n1866), .B0(n1865), .Y(n1874) );
  NAND2X1 U300 ( .A(n1857), .B(n1858), .Y(n1868) );
  OAI31X1 U301 ( .A0(n380), .A1(n379), .A2(n713), .B0(n378), .Y(n413) );
  CLKINVX1 U302 ( .A(curr_time[10]), .Y(n713) );
  NAND2X1 U303 ( .A(n1927), .B(n1929), .Y(n1940) );
  AOI2BB1X2 U304 ( .A0N(n1713), .A1N(n1712), .B0(n1711), .Y(n1721) );
  NOR2X1 U305 ( .A(n880), .B(n879), .Y(n892) );
  OAI31X1 U306 ( .A0(n880), .A1(n879), .A2(n1287), .B0(n878), .Y(n896) );
  OA21X1 U307 ( .A0(n865), .A1(n864), .B0(n863), .Y(n879) );
  OAI31X1 U308 ( .A0(n2220), .A1(n2219), .A2(n2229), .B0(n2218), .Y(n2222) );
  CLKINVX1 U309 ( .A(n2208), .Y(n2220) );
  CLKINVX1 U310 ( .A(n1658), .Y(n1654) );
  OAI211X1 U311 ( .A0(n1332), .A1(n1331), .B0(n690), .C0(n1333), .Y(n2313) );
  NAND2X1 U312 ( .A(n1332), .B(n1331), .Y(n1333) );
  NOR2X1 U313 ( .A(n2318), .B(n2320), .Y(n2319) );
  OAI21X1 U314 ( .A0(n167), .A1(n234), .B0(n2114), .Y(n1373) );
  CLKINVX1 U315 ( .A(n2112), .Y(n2114) );
  CLKINVX1 U316 ( .A(n906), .Y(n916) );
  NAND2X1 U317 ( .A(n2133), .B(n2136), .Y(n2141) );
  NOR2X1 U318 ( .A(n685), .B(n1362), .Y(n1365) );
  CLKINVX1 U319 ( .A(n1208), .Y(n114) );
  NOR2X1 U320 ( .A(n2195), .B(n2204), .Y(n2206) );
  NOR2X1 U321 ( .A(n1636), .B(n1641), .Y(n1648) );
  OAI31X1 U322 ( .A0(n1427), .A1(work_cntr[10]), .A2(n1426), .B0(n1425), .Y(
        n1432) );
  NAND2X1 U323 ( .A(n1416), .B(n1417), .Y(n1427) );
  NOR2X1 U324 ( .A(n1646), .B(n1645), .Y(n1655) );
  CLKINVX1 U325 ( .A(n1949), .Y(n1867) );
  NOR2X1 U326 ( .A(n1565), .B(n1566), .Y(n1588) );
  NAND2X1 U327 ( .A(curr_time[23]), .B(n918), .Y(n305) );
  NOR2X1 U328 ( .A(curr_time[21]), .B(curr_time[22]), .Y(n918) );
  NAND2X1 U329 ( .A(n865), .B(n1771), .Y(n868) );
  OAI31X1 U330 ( .A0(n819), .A1(n818), .A2(n1257), .B0(n817), .Y(n835) );
  OA21X1 U331 ( .A0(n806), .A1(n805), .B0(n804), .Y(n818) );
  NAND2X1 U332 ( .A(n1519), .B(n1582), .Y(n1521) );
  NAND2X1 U333 ( .A(n1549), .B(n1578), .Y(n1557) );
  CLKINVX1 U334 ( .A(n769), .Y(n1780) );
  OAI21X2 U335 ( .A0(n885), .A1(n227), .B0(n756), .Y(n769) );
  NOR2X1 U336 ( .A(n1629), .B(n1628), .Y(n1638) );
  NOR2X1 U337 ( .A(n2292), .B(n257), .Y(n2293) );
  NAND2X1 U338 ( .A(N1233), .B(N1232), .Y(n2292) );
  NOR2X1 U339 ( .A(n2155), .B(n2145), .Y(n2153) );
  NOR2BX1 U340 ( .AN(n2154), .B(n2149), .Y(n2145) );
  AOI2BB2X2 U341 ( .B0(work_cntr[17]), .B1(n1066), .A0N(work_cntr[17]), .A1N(
        n1066), .Y(n1073) );
  NOR2X1 U342 ( .A(n1565), .B(n1587), .Y(n1567) );
  NOR2X1 U343 ( .A(n751), .B(n755), .Y(n753) );
  NAND2X1 U344 ( .A(n2340), .B(n2122), .Y(n2236) );
  NOR2X1 U345 ( .A(n763), .B(n762), .Y(n970) );
  CLKINVX1 U346 ( .A(n1953), .Y(n1908) );
  NOR2BX1 U347 ( .AN(n1810), .B(n1809), .Y(n1818) );
  NOR2X1 U348 ( .A(n1664), .B(n1663), .Y(n1670) );
  NOR2BX1 U349 ( .AN(n2142), .B(n2148), .Y(n2146) );
  NAND2X1 U350 ( .A(n1360), .B(n1359), .Y(n1361) );
  NAND3X1 U351 ( .A(n1010), .B(n1026), .C(n1023), .Y(n1011) );
  AOI31X1 U352 ( .A0(work_cntr[4]), .A1(n2340), .A2(n2119), .B0(
        next_work_cntr[5]), .Y(n2217) );
  NOR2X1 U353 ( .A(n277), .B(n1947), .Y(next_work_cntr[5]) );
  NAND2X1 U354 ( .A(n1683), .B(n1682), .Y(n1688) );
  NOR2X1 U355 ( .A(curr_time[1]), .B(n451), .Y(n437) );
  NAND2X1 U356 ( .A(write_cntr[9]), .B(n766), .Y(n759) );
  OAI31X1 U357 ( .A0(n2246), .A1(n2245), .A2(n2244), .B0(n2243), .Y(n2250) );
  NOR2X1 U358 ( .A(n2251), .B(n2256), .Y(n2244) );
  OAI31X1 U359 ( .A0(n1662), .A1(n1661), .A2(n1660), .B0(n1659), .Y(n1663) );
  NOR2X1 U360 ( .A(n1666), .B(n1665), .Y(n1660) );
  OAI22X1 U361 ( .A0(n1194), .A1(n1193), .B0(n1192), .B1(n1939), .Y(n2326) );
  NOR2X1 U362 ( .A(n1922), .B(n109), .Y(n1194) );
  NOR2X1 U363 ( .A(n2170), .B(n2175), .Y(n2173) );
  AND2X2 U364 ( .A(n2171), .B(n2174), .Y(n2170) );
  NOR2X1 U365 ( .A(n704), .B(n703), .Y(n734) );
  NAND2X1 U366 ( .A(n2209), .B(n2208), .Y(n2226) );
  NAND2BX1 U367 ( .AN(n2202), .B(n2201), .Y(n2208) );
  NAND2BX1 U368 ( .AN(n2201), .B(n2202), .Y(n2209) );
  OAI31X1 U369 ( .A0(n799), .A1(n798), .A2(n1248), .B0(n797), .Y(n811) );
  NAND2X1 U370 ( .A(n261), .B(n193), .Y(n798) );
  OAI31X1 U371 ( .A0(n2252), .A1(n2265), .A2(n2251), .B0(n2264), .Y(n2259) );
  NOR2X1 U372 ( .A(n277), .B(N2063), .Y(n2252) );
  NOR2X1 U373 ( .A(n246), .B(n1317), .Y(n1318) );
  OA21X2 U374 ( .A0(n1969), .A1(n219), .B0(n1626), .Y(n1632) );
  AND2X2 U375 ( .A(n373), .B(n375), .Y(n933) );
  AOI21X1 U376 ( .A0(n249), .A1(n2302), .B0(n2301), .Y(n2306) );
  NOR2BX1 U377 ( .AN(n2129), .B(next_work_cntr[19]), .Y(n2268) );
  OAI31X1 U378 ( .A0(n1724), .A1(n1723), .A2(n1732), .B0(n1722), .Y(n1725) );
  NOR2BX1 U379 ( .AN(n1726), .B(n1729), .Y(n1732) );
  NAND2BX1 U380 ( .AN(n2177), .B(n2176), .Y(n2185) );
  NAND2X1 U381 ( .A(n1582), .B(write_cntr[9]), .Y(n1523) );
  CLKINVX1 U382 ( .A(n1518), .Y(n1582) );
  NOR2X1 U383 ( .A(n177), .B(n1984), .Y(n1994) );
  NAND2X1 U384 ( .A(n1978), .B(n1977), .Y(n1984) );
  AOI2BB2X2 U385 ( .B0(next_work_cntr[9]), .B1(n2123), .A0N(next_work_cntr[9]), 
        .A1N(n2123), .Y(n2194) );
  NAND2X1 U386 ( .A(n2191), .B(n2192), .Y(n2123) );
  NAND3X1 U387 ( .A(n1039), .B(n1026), .C(n1027), .Y(n1028) );
  NOR2X1 U388 ( .A(n2334), .B(n1609), .Y(n1747) );
  INVX3 U389 ( .A(n1772), .Y(n115) );
  NOR2X1 U390 ( .A(n1978), .B(n1977), .Y(n1980) );
  NAND2X2 U391 ( .A(n1672), .B(n214), .Y(n1671) );
  NOR2BX1 U392 ( .AN(n999), .B(n1217), .Y(n1000) );
  NAND2X1 U393 ( .A(n407), .B(n406), .Y(n444) );
  AOI21X1 U394 ( .A0(n214), .A1(n948), .B0(n949), .Y(n1859) );
  NOR2X1 U395 ( .A(n214), .B(n948), .Y(n949) );
  INVXL U396 ( .A(n765), .Y(n116) );
  INVXL U397 ( .A(n116), .Y(n117) );
  NOR2X1 U398 ( .A(n1070), .B(n1069), .Y(n1074) );
  NOR2X1 U399 ( .A(n1067), .B(n177), .Y(n1070) );
  NOR2X1 U400 ( .A(work_cntr[17]), .B(n1982), .Y(n1973) );
  NOR2X1 U401 ( .A(n381), .B(n382), .Y(n412) );
  NOR2BX1 U402 ( .AN(n2097), .B(n2096), .Y(n2099) );
  NOR2X1 U403 ( .A(N2062), .B(N2061), .Y(n2096) );
  OAI21X1 U404 ( .A0(n1385), .A1(n1384), .B0(n1383), .Y(n1391) );
  NAND2X1 U405 ( .A(n1770), .B(n900), .Y(n901) );
  NAND2X1 U406 ( .A(n1326), .B(n1325), .Y(n1329) );
  NOR2X1 U407 ( .A(n1358), .B(n1317), .Y(n1325) );
  NOR2BX1 U408 ( .AN(n1641), .B(n1633), .Y(n1651) );
  NOR2X1 U409 ( .A(n1632), .B(n1630), .Y(n1633) );
  AOI21X1 U410 ( .A0(n2302), .A1(n2297), .B0(n2295), .Y(n2298) );
  NOR2BX1 U411 ( .AN(n1448), .B(n1447), .Y(n1454) );
  NOR2BX1 U412 ( .AN(n1445), .B(n1444), .Y(n1447) );
  OAI21X1 U413 ( .A0(n1504), .A1(n1500), .B0(n187), .Y(n1497) );
  OAI21X1 U414 ( .A0(n1933), .A1(n1932), .B0(n1934), .Y(n1936) );
  NOR2BX1 U415 ( .AN(n1224), .B(n1223), .Y(n1234) );
  OAI21X1 U416 ( .A0(n215), .A1(n1413), .B0(n1410), .Y(n1418) );
  NOR2X1 U417 ( .A(n2194), .B(n2193), .Y(n2205) );
  OAI21X1 U418 ( .A0(n2190), .A1(n2189), .B0(n2188), .Y(n2193) );
  OAI21X1 U419 ( .A0(n265), .A1(n571), .B0(n563), .Y(n521) );
  NOR2BX1 U420 ( .AN(n987), .B(n163), .Y(n988) );
  AND2X2 U421 ( .A(n845), .B(n844), .Y(n848) );
  AOI32X1 U422 ( .A0(n846), .A1(n847), .A2(n845), .B0(n844), .B1(n847), .Y(
        n860) );
  AOI22X1 U423 ( .A0(n2017), .A1(n2016), .B0(n2015), .B1(n2014), .Y(n2021) );
  OAI21X1 U424 ( .A0(n1863), .A1(n1862), .B0(n1861), .Y(n1869) );
  INVXL U425 ( .A(n1887), .Y(n118) );
  INVXL U426 ( .A(n1491), .Y(n119) );
  INVXL U427 ( .A(n1842), .Y(n120) );
  OAI21X1 U428 ( .A0(n1840), .A1(n1844), .B0(n1839), .Y(n1847) );
  INVXL U429 ( .A(n1904), .Y(n121) );
  OAI21X1 U430 ( .A0(n1902), .A1(n1906), .B0(n1901), .Y(n1910) );
  OAI21X1 U431 ( .A0(n1101), .A1(n1108), .B0(n1100), .Y(n1112) );
  NAND3X1 U432 ( .A(write_cntr[1]), .B(write_cntr[0]), .C(write_cntr[2]), .Y(
        n881) );
  NAND2X1 U433 ( .A(n1051), .B(n1048), .Y(n1218) );
  OAI21X1 U434 ( .A0(n1035), .A1(n1034), .B0(n1033), .Y(n1048) );
  NOR2X1 U435 ( .A(N2061), .B(n1498), .Y(n1499) );
  OAI21X1 U436 ( .A0(n167), .A1(n1494), .B0(n1493), .Y(n1498) );
  NOR2X1 U437 ( .A(n1423), .B(n1428), .Y(n1429) );
  OAI21X1 U438 ( .A0(n1422), .A1(n1421), .B0(n1420), .Y(n1428) );
  NOR2X1 U439 ( .A(n277), .B(n1960), .Y(next_work_cntr[13]) );
  OAI211X1 U440 ( .A0(n980), .A1(n256), .B0(n503), .C0(n470), .Y(n501) );
  OAI21X1 U441 ( .A0(n1469), .A1(n1468), .B0(n1467), .Y(n1474) );
  OAI21X1 U442 ( .A0(n1397), .A1(n1396), .B0(n1395), .Y(n1402) );
  INVXL U443 ( .A(n1415), .Y(n122) );
  OAI21X1 U444 ( .A0(n1918), .A1(n1917), .B0(n1916), .Y(n1926) );
  OAI21X1 U445 ( .A0(n1302), .A1(n1301), .B0(n1300), .Y(\intadd_4/B[3] ) );
  AOI22X1 U446 ( .A0(n1188), .A1(n1187), .B0(n1186), .B1(n1185), .Y(n1191) );
  OAI21X1 U447 ( .A0(n1911), .A1(n1183), .B0(n1182), .Y(n1188) );
  OAI22X1 U448 ( .A0(n1145), .A1(n1155), .B0(n1144), .B1(n1143), .Y(n1158) );
  OAI21X1 U449 ( .A0(n1134), .A1(n1133), .B0(n1132), .Y(n1144) );
  OAI22X1 U450 ( .A0(n2020), .A1(n2027), .B0(n2019), .B1(n2018), .Y(n2029) );
  OAI21X1 U451 ( .A0(n2006), .A1(n2014), .B0(n2022), .Y(n2019) );
  NOR2X1 U452 ( .A(n1495), .B(n1499), .Y(n1504) );
  OAI21X1 U453 ( .A0(n1489), .A1(n1493), .B0(n1488), .Y(n1495) );
  NOR2X1 U454 ( .A(n1807), .B(n1806), .Y(n1809) );
  OAI21X1 U455 ( .A0(n1800), .A1(n1804), .B0(n1799), .Y(n1807) );
  OAI211X1 U456 ( .A0(n2106), .A1(n2107), .B0(n2105), .C0(n2104), .Y(n2111) );
  AOI31X1 U457 ( .A0(n1967), .A1(n1966), .A2(n1965), .B0(next_work_cntr[1]), 
        .Y(n2277) );
  OAI21X1 U458 ( .A0(n750), .A1(n1353), .B0(n265), .Y(n2290) );
  BUFX4 U459 ( .A(n1352), .Y(n265) );
  CLKINVX1 U460 ( .A(n512), .Y(n504) );
  NOR2X1 U461 ( .A(read_cntr[1]), .B(n170), .Y(n512) );
  OAI2BB1X2 U462 ( .A0N(n178), .A1N(n945), .B0(n944), .Y(n1948) );
  AOI21X1 U463 ( .A0(n176), .A1(n944), .B0(n947), .Y(n1877) );
  NAND2X1 U464 ( .A(n1969), .B(n219), .Y(n1626) );
  AOI21X1 U465 ( .A0(work_cntr[15]), .A1(n1626), .B0(n1981), .Y(n1629) );
  NAND3X1 U466 ( .A(work_cntr[6]), .B(n1606), .C(n1708), .Y(n944) );
  OAI21X1 U467 ( .A0(n2239), .A1(n2246), .B0(n2238), .Y(n2240) );
  OAI21X1 U468 ( .A0(n1676), .A1(n1669), .B0(n1668), .Y(n1673) );
  INVXL U469 ( .A(n183), .Y(n123) );
  OAI21X1 U470 ( .A0(n1214), .A1(n1213), .B0(n1212), .Y(n1215) );
  NOR2X1 U471 ( .A(work_cntr[10]), .B(n2024), .Y(n2008) );
  OAI21X1 U472 ( .A0(n1816), .A1(n1815), .B0(n1814), .Y(n1823) );
  OAI21X1 U473 ( .A0(n1809), .A1(n1808), .B0(n1951), .Y(n1815) );
  OAI21X1 U474 ( .A0(n1119), .A1(n1118), .B0(n1126), .Y(n1130) );
  OAI21X1 U475 ( .A0(n1447), .A1(n1446), .B0(n176), .Y(n1451) );
  OAI21X1 U476 ( .A0(n1452), .A1(n1451), .B0(n1450), .Y(n1458) );
  NOR2X1 U477 ( .A(work_cntr[13]), .B(n1096), .Y(n1078) );
  OAI21X1 U478 ( .A0(n1267), .A1(n1266), .B0(n1265), .Y(n1270) );
  NAND2BX1 U479 ( .AN(n2127), .B(n2126), .Y(n2128) );
  CLKINVX1 U480 ( .A(next_work_cntr[13]), .Y(n2126) );
  MXI2X2 U481 ( .A(n728), .B(n727), .S0(global_cntr[19]), .Y(next_glb_cntr[19]) );
  OAI21X1 U482 ( .A0(n1524), .A1(n1536), .B0(n1523), .Y(n1525) );
  NOR2X1 U483 ( .A(write_cntr[9]), .B(n1582), .Y(n1524) );
  NAND2X1 U484 ( .A(n868), .B(n866), .Y(n874) );
  OAI22X1 U485 ( .A0(n1027), .A1(n853), .B0(n852), .B1(n851), .Y(n866) );
  NOR2X4 U486 ( .A(n1368), .B(n2330), .Y(n645) );
  NAND2XL U487 ( .A(N473), .B(\DP_OP_665J1_134_4923/I2 ), .Y(
        \DP_OP_665J1_134_4923/n111 ) );
  OAI21X1 U488 ( .A0(N2061), .A1(n1738), .B0(n1742), .Y(n1754) );
  OAI22X1 U489 ( .A0(n2096), .A1(n1737), .B0(n1736), .B1(n1735), .Y(n1738) );
  NOR2X2 U490 ( .A(n751), .B(n721), .Y(n1764) );
  NAND2X1 U491 ( .A(n2216), .B(n2215), .Y(n2225) );
  OAI22X1 U492 ( .A0(n2214), .A1(n2213), .B0(n2212), .B1(n2211), .Y(n2215) );
  OAI22X1 U493 ( .A0(n1939), .A1(n1750), .B0(n1741), .B1(n1754), .Y(
        expand_sel[1]) );
  NAND2X1 U494 ( .A(n1609), .B(n1608), .Y(n1750) );
  NOR3X1 U495 ( .A(n1606), .B(n1605), .C(n2334), .Y(n1608) );
  CLKINVX1 U496 ( .A(n2087), .Y(n2092) );
  OAI22X1 U497 ( .A0(work_cntr[4]), .A1(n2076), .B0(n180), .B1(n2077), .Y(
        n2087) );
  AOI2BB1X2 U498 ( .A0N(work_cntr[4]), .A1N(n1606), .B0(n946), .Y(n1953) );
  NOR2X1 U499 ( .A(n180), .B(n2119), .Y(n946) );
  AOI31X1 U500 ( .A0(n2164), .A1(n2163), .A2(n2162), .B0(n2161), .Y(n2167) );
  CLKINVX1 U501 ( .A(n2058), .Y(n1687) );
  OAI21X1 U502 ( .A0(n1667), .A1(n1663), .B0(n1664), .Y(n1678) );
  NOR3BX1 U503 ( .AN(n1664), .B(n1679), .C(n1665), .Y(n1667) );
  OAI21X1 U504 ( .A0(n996), .A1(n1008), .B0(n995), .Y(n997) );
  OAI21X1 U505 ( .A0(n988), .A1(N585), .B0(n1356), .Y(n1354) );
  OAI31X4 U506 ( .A0(n858), .A1(n857), .A2(n1274), .B0(n856), .Y(n872) );
  AOI2BB2X2 U507 ( .B0(n998), .B1(n997), .A0N(n998), .A1N(n997), .Y(n1012) );
  OAI22X2 U508 ( .A0(n1779), .A1(n1230), .B0(n961), .B1(next_cr_x[6]), .Y(n998) );
  NAND2X1 U509 ( .A(n1720), .B(n180), .Y(n1728) );
  OAI31X1 U510 ( .A0(n1719), .A1(n1718), .A2(n1717), .B0(n1716), .Y(n1720) );
  NOR2X1 U511 ( .A(n2199), .B(n2205), .Y(n2195) );
  NOR3X1 U512 ( .A(n2194), .B(n2204), .C(n2197), .Y(n2199) );
  NOR3BX1 U513 ( .AN(n1694), .B(n1707), .C(n1689), .Y(n1701) );
  OAI21X2 U514 ( .A0(n1687), .A1(n176), .B0(n2041), .Y(n1694) );
  NOR2X1 U515 ( .A(n2250), .B(n2249), .Y(n2260) );
  NOR3BX1 U516 ( .AN(n2143), .B(n2155), .C(n2147), .Y(n2149) );
  AOI32X1 U517 ( .A0(n2262), .A1(n2254), .A2(n2253), .B0(n2259), .B1(n2254), 
        .Y(n2263) );
  OAI31X1 U518 ( .A0(n838), .A1(n1264), .A2(n837), .B0(n836), .Y(n846) );
  NOR2X1 U519 ( .A(n215), .B(n951), .Y(n952) );
  OAI21X1 U520 ( .A0(n1462), .A1(n1454), .B0(n178), .Y(n1459) );
  OA21X2 U521 ( .A0(n178), .A1(n1461), .B0(n1459), .Y(n1469) );
  OAI31X4 U522 ( .A0(n1037), .A1(\intadd_3/A[0] ), .A2(n1771), .B0(n1036), .Y(
        n1038) );
  AOI2BB2X2 U523 ( .B0(n1010), .B1(n1009), .A0N(n1010), .A1N(n1009), .Y(n1030)
         );
  NAND2X1 U524 ( .A(n938), .B(n713), .Y(n937) );
  MXI2X1 U525 ( .A(n932), .B(curr_time[11]), .S0(n933), .Y(n938) );
  NOR4X1 U526 ( .A(n698), .B(n697), .C(n696), .D(n695), .Y(n735) );
  AOI211X1 U527 ( .A0(n2324), .A1(n2323), .B0(n2322), .C0(n2325), .Y(n2333) );
  OA22X2 U528 ( .A0(n885), .A1(n211), .B0(n270), .B1(n754), .Y(n175) );
  NOR2X1 U529 ( .A(n321), .B(n320), .Y(n375) );
  NOR2X1 U530 ( .A(n369), .B(n368), .Y(n681) );
  NOR2X1 U531 ( .A(n966), .B(n967), .Y(n965) );
  NOR2X1 U532 ( .A(n1168), .B(n1167), .Y(n1174) );
  AOI21X1 U533 ( .A0(n1174), .A1(n1177), .B0(n1169), .Y(n1181) );
  NOR2X1 U534 ( .A(n210), .B(n775), .Y(n780) );
  NOR2X1 U535 ( .A(n1099), .B(n1107), .Y(n1115) );
  AOI21X1 U536 ( .A0(n1107), .A1(n1106), .B0(n1115), .Y(n1110) );
  AOI2BB2X2 U537 ( .B0(next_work_cntr[11]), .B1(n2125), .A0N(
        next_work_cntr[11]), .A1N(n2125), .Y(n2176) );
  NOR2BX1 U538 ( .AN(n2124), .B(next_work_cntr[10]), .Y(n2125) );
  NOR2X1 U539 ( .A(n819), .B(n818), .Y(n824) );
  NAND3X1 U540 ( .A(write_cntr[9]), .B(write_cntr[11]), .C(write_cntr[10]), 
        .Y(n1519) );
  OAI211X1 U541 ( .A0(write_cntr[11]), .A1(n757), .B0(n755), .C0(n783), .Y(
        n756) );
  NOR2X1 U542 ( .A(n1985), .B(n1994), .Y(n1991) );
  NOR2X1 U543 ( .A(n412), .B(n411), .Y(n457) );
  NOR2X1 U544 ( .A(n799), .B(n798), .Y(n802) );
  NOR2X1 U545 ( .A(n792), .B(n793), .Y(n799) );
  AOI21X1 U546 ( .A0(n171), .A1(n745), .B0(n691), .Y(n1060) );
  AOI2BB2X2 U547 ( .B0(n2165), .B1(next_work_cntr[12]), .A0N(n2165), .A1N(
        next_work_cntr[12]), .Y(n2166) );
  NAND2BX1 U548 ( .AN(next_work_cntr[12]), .B(n2165), .Y(n2127) );
  NOR2BX1 U549 ( .AN(n2125), .B(next_work_cntr[11]), .Y(n2165) );
  NOR2X1 U550 ( .A(n1060), .B(n1059), .Y(n1065) );
  AOI21X1 U551 ( .A0(n1140), .A1(n1139), .B0(n1146), .Y(n1142) );
  NOR2X1 U552 ( .A(n1131), .B(n1140), .Y(n1146) );
  OAI22X1 U553 ( .A0(n1623), .A1(n1622), .B0(n1621), .B1(n1620), .Y(n1628) );
  CLKINVX1 U554 ( .A(n2257), .Y(n2251) );
  OAI2BB2X1 U555 ( .B0(n2236), .B1(n2235), .A0N(n2236), .A1N(n2235), .Y(n2257)
         );
  OAI21X1 U556 ( .A0(n1973), .A1(n177), .B0(n1971), .Y(n1622) );
  OAI21X1 U557 ( .A0(n2221), .A1(n2222), .B0(n2223), .Y(n2237) );
  NAND2X1 U558 ( .A(n2237), .B(n2238), .Y(n2245) );
  OAI21X1 U559 ( .A0(n916), .A1(n915), .B0(n914), .Y(n1204) );
  AOI221X4 U560 ( .A0(n1206), .A1(n1205), .B0(n1204), .B1(n1205), .C0(n1213), 
        .Y(n1207) );
  AOI2BB2X2 U561 ( .B0(n1199), .B1(n1198), .A0N(n1204), .A1N(n1197), .Y(n1209)
         );
  OAI21X1 U562 ( .A0(n408), .A1(n409), .B0(n444), .Y(n454) );
  OAI21X1 U563 ( .A0(work_cntr[19]), .A1(n1959), .B0(n1786), .Y(n1792) );
  OAI31X1 U564 ( .A0(n1794), .A1(n1793), .A2(n1792), .B0(n1791), .Y(n1802) );
  OAI21X1 U565 ( .A0(n222), .A1(n1417), .B0(n1421), .Y(n1426) );
  OAI21X1 U566 ( .A0(n2057), .A1(n178), .B0(n2058), .Y(n1705) );
  OAI21X1 U567 ( .A0(n168), .A1(n1465), .B0(n1468), .Y(n1472) );
  CLKINVX1 U568 ( .A(n1147), .Y(n1133) );
  AOI2BB2X2 U569 ( .B0(n1142), .B1(n1141), .A0N(n1142), .A1N(n1147), .Y(n1154)
         );
  OAI2BB2X1 U570 ( .B0(n1705), .B1(n1709), .A0N(n1705), .A1N(n1709), .Y(n1724)
         );
  OAI2BB2X1 U571 ( .B0(work_cntr[8]), .B1(n1135), .A0N(work_cntr[8]), .A1N(
        n1135), .Y(n1147) );
  OAI221X1 U572 ( .A0(n1087), .A1(n1090), .B0(n1083), .B1(n1090), .C0(n1082), 
        .Y(n1086) );
  OAI21X1 U573 ( .A0(n1076), .A1(n181), .B0(n1075), .Y(n1087) );
  NOR2BX1 U574 ( .AN(n1082), .B(n1087), .Y(n1091) );
  OAI21X1 U575 ( .A0(n219), .A1(n1393), .B0(n1396), .Y(n1400) );
  OAI21X1 U576 ( .A0(n1122), .A1(n1121), .B0(n1120), .Y(n1125) );
  OAI21X1 U577 ( .A0(n265), .A1(n2310), .B0(n2311), .Y(n629) );
  OAI2BB2X1 U578 ( .B0(n1110), .B1(n1116), .A0N(n1110), .A1N(n1109), .Y(n1122)
         );
  OAI21X1 U579 ( .A0(n1078), .A1(n219), .B0(n1077), .Y(n1088) );
  OAI2BB2X1 U580 ( .B0(n1442), .B1(n1438), .A0N(n1442), .A1N(n1438), .Y(n1444)
         );
  OAI21X1 U581 ( .A0(n214), .A1(n1436), .B0(n1434), .Y(n1438) );
  NOR3X1 U582 ( .A(n1629), .B(n1631), .C(n1616), .Y(n1624) );
  OAI2BB2X1 U583 ( .B0(next_work_cntr[10]), .B1(n2124), .A0N(
        next_work_cntr[10]), .A1N(n2124), .Y(n2183) );
  OAI22X1 U584 ( .A0(n1530), .A1(n1529), .B0(n1531), .B1(n1533), .Y(n1546) );
  OAI22X1 U585 ( .A0(n1022), .A1(n1021), .B0(n1032), .B1(n1020), .Y(n1049) );
  OAI31X1 U586 ( .A0(n1596), .A1(n1574), .A2(n1597), .B0(n1586), .Y(n1583) );
  OAI22X1 U587 ( .A0(n717), .A1(n1576), .B0(n1573), .B1(n1572), .Y(n1586) );
  OAI21X1 U588 ( .A0(n1264), .A1(n1263), .B0(n1262), .Y(n1272) );
  NOR2X1 U589 ( .A(n994), .B(n822), .Y(n819) );
  OAI22X1 U590 ( .A0(n1252), .A1(n1779), .B0(n1251), .B1(n961), .Y(n822) );
  NAND2X1 U591 ( .A(n901), .B(n904), .Y(n895) );
  OAI22X1 U592 ( .A0(n1040), .A1(n889), .B0(n888), .B1(n887), .Y(n904) );
  OAI31X1 U593 ( .A0(n913), .A1(n912), .A2(n911), .B0(n910), .Y(n1214) );
  NAND2BX1 U594 ( .AN(n913), .B(n912), .Y(n915) );
  OAI22X1 U595 ( .A0(n903), .A1(n901), .B0(n900), .B1(n899), .Y(n912) );
  OAI22X1 U596 ( .A0(n1983), .A1(n182), .B0(n1982), .B1(n2077), .Y(n1993) );
  CLKINVX1 U597 ( .A(n898), .Y(n1770) );
  OAI22X1 U598 ( .A0(n225), .A1(n885), .B0(n270), .B1(n883), .Y(n898) );
  AOI32X1 U599 ( .A0(n810), .A1(n809), .A2(n808), .B0(n807), .B1(n809), .Y(
        n825) );
  OAI21X1 U600 ( .A0(n802), .A1(n801), .B0(n800), .Y(n810) );
  OAI22X1 U601 ( .A0(work_cntr[10]), .A1(n1610), .B0(n183), .B1(n1671), .Y(
        n1674) );
  AOI2BB2X2 U602 ( .B0(n2182), .B1(n2184), .A0N(n2182), .A1N(n2184), .Y(n2204)
         );
  NOR2X1 U603 ( .A(n2184), .B(n2183), .Y(n2196) );
  OAI31X4 U604 ( .A0(n2187), .A1(n2181), .A2(n2180), .B0(n2179), .Y(n2184) );
  OA21X2 U605 ( .A0(n419), .A1(n418), .B0(n421), .Y(n451) );
  OAI21X1 U606 ( .A0(n896), .A1(n895), .B0(n894), .Y(n911) );
  OAI21X1 U607 ( .A0(n892), .A1(n891), .B0(n890), .Y(n897) );
  OAI31X1 U608 ( .A0(n871), .A1(n870), .A2(n1285), .B0(n869), .Y(n891) );
  OAI31X1 U609 ( .A0(n1287), .A1(n1298), .A2(n1299), .B0(n1286), .Y(
        \intadd_4/A[2] ) );
  OAI31X4 U610 ( .A0(n1285), .A1(n1284), .A2(n1283), .B0(n1282), .Y(n1299) );
  NAND2X1 U611 ( .A(n833), .B(n829), .Y(n837) );
  NAND2BX1 U612 ( .AN(n1695), .B(n1694), .Y(n1706) );
  AOI2BB2X2 U613 ( .B0(n1694), .B1(n1695), .A0N(n1694), .A1N(n1695), .Y(n1717)
         );
  OAI31X4 U614 ( .A0(n1701), .A1(n1693), .A2(n1692), .B0(n1691), .Y(n1695) );
  CLKINVX1 U615 ( .A(n849), .Y(n125) );
  CLKINVX1 U616 ( .A(n125), .Y(n126) );
  CLKINVX1 U617 ( .A(n1378), .Y(n127) );
  CLKINVX1 U618 ( .A(n127), .Y(n128) );
  CLKINVX1 U619 ( .A(n1747), .Y(n1741) );
  XOR2X1 U620 ( .A(n981), .B(n271), .Y(n1328) );
  CLKINVX1 U621 ( .A(n671), .Y(\im_a[1]_BAR ) );
  CLKINVX1 U622 ( .A(n673), .Y(\im_a[2]_BAR ) );
  CLKINVX1 U623 ( .A(n675), .Y(\im_a[17]_BAR ) );
  OAI2BB2X1 U624 ( .B0(next_work_cntr[18]), .B1(n2130), .A0N(
        next_work_cntr[18]), .A1N(n2130), .Y(n2138) );
  NOR2X1 U625 ( .A(n2130), .B(next_work_cntr[18]), .Y(n2129) );
  NOR2X2 U626 ( .A(n277), .B(n1965), .Y(next_work_cntr[18]) );
  NOR3X2 U627 ( .A(n460), .B(n459), .C(n458), .Y(\DP_OP_251J1_126_494/I2 ) );
  CLKINVX1 U628 ( .A(n404), .Y(n460) );
  CLKINVX1 U629 ( .A(n1511), .Y(n572) );
  NOR2X2 U630 ( .A(n691), .B(n1370), .Y(n1511) );
  OAI2BB2X1 U631 ( .B0(curr_time[4]), .B1(\s_1[3] ), .A0N(curr_time[4]), .A1N(
        \s_1[3] ), .Y(n943) );
  NAND2X1 U632 ( .A(n323), .B(n387), .Y(\s_1[3] ) );
  OAI21X1 U633 ( .A0(n1172), .A1(n1171), .B0(n1173), .Y(n1178) );
  NAND2X1 U634 ( .A(n1168), .B(n1171), .Y(n1173) );
  OAI21X2 U635 ( .A0(n1157), .A1(n168), .B0(n1156), .Y(n1171) );
  OAI31X1 U636 ( .A0(n814), .A1(n1251), .A2(n813), .B0(n812), .Y(n816) );
  NAND2X1 U637 ( .A(n808), .B(n807), .Y(n813) );
  OAI21X2 U638 ( .A0(n2333), .A1(n2336), .B0(n2335), .Y(so_mux_sel[0]) );
  CLKINVX1 U639 ( .A(curr_time[18]), .Y(n711) );
  OAI21X1 U640 ( .A0(n1612), .A1(n215), .B0(n1634), .Y(n1658) );
  NOR2X2 U641 ( .A(work_cntr[13]), .B(n1634), .Y(n1969) );
  NAND2X1 U642 ( .A(n1612), .B(n215), .Y(n1634) );
  OAI2BB2X1 U643 ( .B0(curr_time[20]), .B1(h_1[3]), .A0N(curr_time[20]), .A1N(
        h_1[3]), .Y(n924) );
  NAND2X1 U644 ( .A(n301), .B(n305), .Y(h_1[3]) );
  OAI21X2 U645 ( .A0(n1073), .A1(n1072), .B0(n1071), .Y(n1080) );
  OAI21X1 U646 ( .A0(work_cntr[19]), .A1(n1070), .B0(n1069), .Y(n1072) );
  OAI21X2 U647 ( .A0(\intadd_3/SUM[4] ), .A1(n1353), .B0(n186), .Y(n621) );
  NOR3X2 U648 ( .A(n403), .B(n1768), .C(n1767), .Y(n459) );
  NAND2X1 U649 ( .A(n458), .B(n403), .Y(n440) );
  NAND2X1 U650 ( .A(n1599), .B(n1600), .Y(n403) );
  NAND2X1 U651 ( .A(n179), .B(n1725), .Y(n1745) );
  NAND2X1 U652 ( .A(write_addr[8]), .B(n1361), .Y(n1370) );
  NOR3X1 U653 ( .A(write_addr[8]), .B(n685), .C(n1373), .Y(n1364) );
  OAI21X1 U654 ( .A0(n2075), .A1(n2082), .B0(n2090), .Y(n2088) );
  AOI22X1 U655 ( .A0(n2085), .A1(n2084), .B0(n2083), .B1(n2082), .Y(n2089) );
  OAI22X2 U656 ( .A0(n2061), .A1(n168), .B0(n2060), .B1(n2077), .Y(n2082) );
  OAI21X1 U657 ( .A0(n2056), .A1(n2066), .B0(n2074), .Y(n2071) );
  AOI22X1 U658 ( .A0(n2069), .A1(n2068), .B0(n2067), .B1(n2066), .Y(n2073) );
  OAI22X2 U659 ( .A0(n2042), .A1(n176), .B0(n2041), .B1(n2077), .Y(n2066) );
  OAI21X1 U660 ( .A0(n2039), .A1(n2047), .B0(n2055), .Y(n2052) );
  AOI22X1 U661 ( .A0(n2050), .A1(n2049), .B0(n2048), .B1(n2047), .Y(n2054) );
  OAI21X2 U662 ( .A0(n2025), .A1(n214), .B0(n2024), .Y(n2047) );
  OAI21X1 U663 ( .A0(n2023), .A1(n2030), .B0(n2038), .Y(n2035) );
  AOI22X1 U664 ( .A0(n2033), .A1(n2032), .B0(n2031), .B1(n2030), .Y(n2037) );
  OAI21X2 U665 ( .A0(n2008), .A1(n222), .B0(n2007), .Y(n2030) );
  NAND2X2 U666 ( .A(n2331), .B(n1739), .Y(n1934) );
  NAND2X1 U667 ( .A(N2062), .B(n1739), .Y(n2323) );
  NOR2X1 U668 ( .A(N2062), .B(n1739), .Y(n1751) );
  NAND2X1 U669 ( .A(n187), .B(n234), .Y(n1739) );
  NOR2X2 U670 ( .A(n277), .B(n1959), .Y(next_work_cntr[17]) );
  AOI211X4 U671 ( .A0(n192), .A1(n689), .B0(n1309), .C0(n352), .Y(n596) );
  OAI22X2 U672 ( .A0(n2059), .A1(n178), .B0(n2058), .B1(n2077), .Y(n2079) );
  NAND2X1 U673 ( .A(n178), .B(n2057), .Y(n2058) );
  OAI21X1 U674 ( .A0(n2064), .A1(n2063), .B0(n2062), .Y(n2067) );
  OAI22X1 U675 ( .A0(n2053), .A1(n2063), .B0(n2052), .B1(n2051), .Y(n2065) );
  OAI2BB2X2 U676 ( .B0(n2040), .B1(n226), .A0N(n2040), .A1N(n226), .Y(n2063)
         );
  OAI2BB2X2 U677 ( .B0(work_cntr[10]), .B1(n2024), .A0N(work_cntr[10]), .A1N(
        n2024), .Y(n2044) );
  NAND2X1 U678 ( .A(n2025), .B(n214), .Y(n2024) );
  OAI2BB2X2 U679 ( .B0(work_cntr[12]), .B1(n2007), .A0N(work_cntr[12]), .A1N(
        n2007), .Y(n2027) );
  NAND2X1 U680 ( .A(n2008), .B(n222), .Y(n2007) );
  AOI2BB2X2 U681 ( .B0(n1315), .B1(write_addr[16]), .A0N(n1315), .A1N(
        write_addr[16]), .Y(n1326) );
  AOI21X1 U682 ( .A0(n247), .A1(n1316), .B0(n1315), .Y(n1320) );
  NOR2X2 U683 ( .A(n1358), .B(n1310), .Y(n1315) );
  OAI2BB2X1 U684 ( .B0(n1196), .B1(\next_cr_y[0] ), .A0N(n1196), .A1N(
        \next_cr_y[0] ), .Y(n1054) );
  OAI22X2 U685 ( .A0(write_cntr[0]), .A1(n270), .B0(n185), .B1(n885), .Y(n1196) );
  CLKINVX1 U686 ( .A(n365), .Y(n682) );
  NOR2X2 U687 ( .A(n355), .B(n354), .Y(n586) );
  NAND2X1 U688 ( .A(n1535), .B(n1579), .Y(n1541) );
  NAND2X1 U689 ( .A(n1609), .B(n2076), .Y(n2112) );
  NOR2X2 U690 ( .A(n1971), .B(work_cntr[19]), .Y(n1609) );
  OAI21X2 U691 ( .A0(n1102), .A1(n215), .B0(n1096), .Y(n1108) );
  NAND2BX1 U692 ( .AN(n1634), .B(n1163), .Y(n1096) );
  ADDFX2 U693 ( .A(n167), .B(n1743), .CI(n1742), .CO(n1760), .S(n1756) );
  NAND2X1 U694 ( .A(n1636), .B(n1635), .Y(n1661) );
  INVXL U695 ( .A(n1528), .Y(n129) );
  CLKINVX1 U696 ( .A(n129), .Y(n130) );
  OAI2BB2X2 U697 ( .B0(n213), .B1(n1982), .A0N(n213), .A1N(n1982), .Y(n1618)
         );
  NAND2X2 U698 ( .A(n1981), .B(n182), .Y(n1982) );
  OAI2BB2X2 U699 ( .B0(n1684), .B1(n1683), .A0N(n1684), .A1N(n1683), .Y(n1700)
         );
  AOI31X4 U700 ( .A0(n1679), .A1(n1678), .A2(n1677), .B0(n1676), .Y(n1683) );
  NOR2X2 U701 ( .A(n277), .B(n1946), .Y(next_work_cntr[10]) );
  OA21X2 U702 ( .A0(n1946), .A1(n1854), .B0(n1848), .Y(n1863) );
  CLKINVX1 U703 ( .A(n1851), .Y(n1946) );
  CLKINVX1 U704 ( .A(n1040), .Y(n1774) );
  CLKINVX1 U705 ( .A(n1337), .Y(n131) );
  NAND2X1 U706 ( .A(n2340), .B(n167), .Y(n2262) );
  CLKINVX1 U707 ( .A(n1338), .Y(n132) );
  OAI22X2 U708 ( .A0(n1002), .A1(n1217), .B0(n1778), .B1(n1237), .Y(n1026) );
  CLKINVX1 U709 ( .A(n1778), .Y(n1002) );
  OAI21X1 U710 ( .A0(n1330), .A1(n165), .B0(n2340), .Y(n1245) );
  NOR3X1 U711 ( .A(n231), .B(n1330), .C(n1329), .Y(n1331) );
  CLKINVX1 U712 ( .A(n1306), .Y(n1330) );
  NAND2X1 U713 ( .A(n1564), .B(n1601), .Y(n1570) );
  NOR2X2 U714 ( .A(n1601), .B(write_cntr[5]), .Y(n1592) );
  OAI21X2 U715 ( .A0(n1989), .A1(n221), .B0(n1988), .Y(n2014) );
  NAND2X1 U716 ( .A(n1969), .B(n2076), .Y(n1988) );
  NOR2X1 U717 ( .A(read_cntr[0]), .B(read_cntr[1]), .Y(n684) );
  OAI211X1 U718 ( .A0(read_cntr[0]), .A1(n1363), .B0(n514), .C0(n513), .Y(n515) );
  OAI21X1 U719 ( .A0(read_cntr[0]), .A1(n233), .B0(n504), .Y(n658) );
  OAI2BB2X1 U720 ( .B0(work_cntr[10]), .B1(n1127), .A0N(work_cntr[10]), .A1N(
        n1127), .Y(n1123) );
  AOI21X1 U721 ( .A0(work_cntr[9]), .A1(n1128), .B0(n1127), .Y(n1140) );
  NOR2X2 U722 ( .A(n1671), .B(n1164), .Y(n1127) );
  OAI31X1 U723 ( .A0(n771), .A1(n1247), .A2(n790), .B0(n789), .Y(n795) );
  NOR2BX1 U724 ( .AN(n771), .B(n790), .Y(n784) );
  NAND2X1 U725 ( .A(n771), .B(n761), .Y(n770) );
  NAND2X1 U726 ( .A(n771), .B(n770), .Y(n968) );
  CLKINVX1 U727 ( .A(n174), .Y(n771) );
  OAI21X2 U728 ( .A0(n2103), .A1(n2102), .B0(n2101), .Y(n2107) );
  OAI21X2 U729 ( .A0(n2097), .A1(n179), .B0(n2077), .Y(n2102) );
  NAND2X1 U730 ( .A(write_cntr[11]), .B(n757), .Y(n755) );
  NOR2X1 U731 ( .A(n107), .B(n759), .Y(n757) );
  AND2X2 U732 ( .A(n1769), .B(n909), .Y(n913) );
  NOR2BX1 U733 ( .AN(n1769), .B(n1240), .Y(n908) );
  AOI21X2 U734 ( .A0(n773), .A1(write_cntr[1]), .B0(n772), .Y(n1769) );
  NOR2X1 U735 ( .A(n1230), .B(n1229), .Y(n1238) );
  NOR2BX1 U736 ( .AN(n1011), .B(n1229), .Y(n1007) );
  OAI22X2 U737 ( .A0(n1023), .A1(n1229), .B0(n1776), .B1(n1231), .Y(n1039) );
  NOR2X1 U738 ( .A(n1229), .B(n1215), .Y(n1221) );
  CLKINVX1 U739 ( .A(n1231), .Y(n1229) );
  NAND3X1 U740 ( .A(write_cntr[6]), .B(n1556), .C(n1569), .Y(n1549) );
  AND2X2 U741 ( .A(n1578), .B(write_cntr[6]), .Y(n1565) );
  OAI21X1 U742 ( .A0(work_cntr[18]), .A1(n956), .B0(n1785), .Y(n1965) );
  OAI2BB2X1 U743 ( .B0(work_cntr[19]), .B1(n1785), .A0N(n1784), .A1N(n1783), 
        .Y(n1789) );
  NAND2X1 U744 ( .A(work_cntr[18]), .B(n956), .Y(n1785) );
  CLKINVX1 U745 ( .A(n649), .Y(n592) );
  NOR2X2 U746 ( .A(n277), .B(n1952), .Y(next_work_cntr[12]) );
  OAI21X1 U747 ( .A0(n1952), .A1(n1836), .B0(n1832), .Y(n1834) );
  CLKINVX1 U748 ( .A(n1829), .Y(n1952) );
  AND3X2 U749 ( .A(state[0]), .B(n28), .C(n205), .Y(n171) );
  OA22X1 U750 ( .A0(n172), .A1(n1059), .B0(state[0]), .B1(n743), .Y(n744) );
  OR2X1 U751 ( .A(state[0]), .B(curr_photo_size[0]), .Y(n325) );
  NOR3X2 U752 ( .A(n123), .B(work_cntr[11]), .C(n1671), .Y(n1612) );
  CLKINVX1 U753 ( .A(n1308), .Y(n690) );
  OAI21X2 U754 ( .A0(work_cntr[13]), .A1(n952), .B0(n953), .Y(n1960) );
  NAND2X2 U755 ( .A(work_cntr[13]), .B(n952), .Y(n953) );
  NAND3X2 U756 ( .A(n467), .B(n466), .C(n465), .Y(\DP_OP_251J1_126_494/I3 ) );
  NAND2X1 U757 ( .A(n459), .B(n1601), .Y(n465) );
  NOR4X1 U758 ( .A(n464), .B(n463), .C(n462), .D(n461), .Y(n467) );
  OAI22X1 U759 ( .A0(n769), .A1(n1247), .B0(n1780), .B1(n784), .Y(n793) );
  OAI31X1 U760 ( .A0(n788), .A1(n787), .A2(n1247), .B0(n786), .Y(n801) );
  AND2X2 U761 ( .A(n1247), .B(n1249), .Y(n184) );
  CLKINVX1 U762 ( .A(n784), .Y(n1247) );
  NOR2X2 U763 ( .A(n2057), .B(n1708), .Y(n2122) );
  NOR2X1 U764 ( .A(n168), .B(n180), .Y(n1708) );
  NOR2X1 U765 ( .A(work_cntr[16]), .B(n1377), .Y(n1381) );
  OAI2BB2X1 U766 ( .B0(work_cntr[16]), .B1(n128), .A0N(work_cntr[16]), .A1N(
        n128), .Y(n1385) );
  AOI221X1 U767 ( .A0(work_cntr[16]), .A1(n1390), .B0(n1380), .B1(n1390), .C0(
        n1379), .Y(n1388) );
  NOR2X2 U768 ( .A(n1075), .B(work_cntr[16]), .Y(n1066) );
  NOR2X1 U769 ( .A(work_cntr[8]), .B(n2041), .Y(n1672) );
  NOR2X2 U770 ( .A(n2041), .B(n1164), .Y(n1135) );
  NOR3X1 U771 ( .A(work_cntr[8]), .B(n2041), .C(n2077), .Y(n2025) );
  AOI21X1 U772 ( .A0(work_cntr[8]), .A1(n2041), .B0(n1672), .Y(n1696) );
  NOR2X1 U773 ( .A(n2041), .B(n2077), .Y(n2040) );
  NAND2X2 U774 ( .A(n1687), .B(n176), .Y(n2041) );
  CLKINVX1 U775 ( .A(n1251), .Y(n1252) );
  NOR2X2 U776 ( .A(n803), .B(n810), .Y(n1251) );
  CLKINVX1 U777 ( .A(n1237), .Y(n1217) );
  NAND2X2 U778 ( .A(n1004), .B(n1003), .Y(n1237) );
  CLKINVX1 U779 ( .A(n115), .Y(n994) );
  OAI22X2 U780 ( .A0(n115), .A1(next_cr_x[5]), .B0(n994), .B1(n1223), .Y(n1010) );
  CLKINVX1 U781 ( .A(en_so), .Y(n663) );
  NAND2X4 U782 ( .A(en_so), .B(state[0]), .Y(n2334) );
  NAND2X4 U783 ( .A(n2328), .B(n742), .Y(en_so) );
  AOI211X4 U784 ( .A0(n348), .A1(N579), .B0(n1202), .C0(n337), .Y(n640) );
  NOR2X1 U785 ( .A(n1934), .B(n277), .Y(next_work_cntr[1]) );
  INVX3 U786 ( .A(n266), .Y(n661) );
  OAI21X1 U787 ( .A0(work_cntr[8]), .A1(n1438), .B0(n1440), .Y(n1441) );
  AOI21X1 U788 ( .A0(n1441), .A1(n1439), .B0(work_cntr[8]), .Y(n1442) );
  NAND2X1 U789 ( .A(n2340), .B(n1867), .Y(n2192) );
  NAND2X1 U790 ( .A(n180), .B(n2340), .Y(n2248) );
  OAI21X1 U791 ( .A0(n179), .A1(n1486), .B0(n1482), .Y(n1484) );
  INVX3 U792 ( .A(n563), .Y(n568) );
  AOI2BB1X4 U793 ( .A0N(n516), .A1N(n1369), .B0(n515), .Y(n563) );
  NAND2X1 U794 ( .A(n1027), .B(n1224), .Y(n1036) );
  OAI21X1 U795 ( .A0(n1224), .A1(n1027), .B0(n1036), .Y(n1042) );
  NAND2X2 U796 ( .A(n1033), .B(n1032), .Y(n1224) );
  INVX16 U797 ( .A(n6), .Y(cr_a[2]) );
  INVX16 U798 ( .A(n5), .Y(cr_a[1]) );
  NAND2X1 U799 ( .A(N2062), .B(N2061), .Y(n2097) );
  INVX16 U800 ( .A(n3), .Y(cr_a[0]) );
  CLKINVX1 U801 ( .A(n2346), .Y(n136) );
  INVX16 U802 ( .A(n136), .Y(cr_a[3]) );
  CLKINVX1 U803 ( .A(n2345), .Y(n138) );
  INVX16 U804 ( .A(n138), .Y(cr_a[4]) );
  CLKINVX1 U805 ( .A(n2344), .Y(n140) );
  INVX16 U806 ( .A(n140), .Y(cr_a[5]) );
  CLKINVX1 U807 ( .A(n2343), .Y(n142) );
  INVX16 U808 ( .A(n142), .Y(cr_a[6]) );
  CLKINVX1 U809 ( .A(n2342), .Y(n144) );
  INVX16 U810 ( .A(n144), .Y(cr_a[7]) );
  INVX16 U811 ( .A(n7), .Y(cr_a[8]) );
  INVX16 U812 ( .A(n2341), .Y(im_wen_n) );
  INVX3 U813 ( .A(n254), .Y(n268) );
  NAND2X1 U814 ( .A(n663), .B(n276), .Y(n254) );
  NAND2BX1 U815 ( .AN(n978), .B(n977), .Y(n980) );
  NOR2X1 U816 ( .A(n189), .B(n974), .Y(n978) );
  NOR2X1 U817 ( .A(n2297), .B(n2296), .Y(n2300) );
  NAND2X1 U818 ( .A(cr_read_cntr[3]), .B(n2294), .Y(n2296) );
  NAND2BX1 U819 ( .AN(n1462), .B(n1461), .Y(n1466) );
  NOR2X1 U820 ( .A(n1453), .B(n1458), .Y(n1462) );
  NAND2BX1 U821 ( .AN(n1824), .B(n1826), .Y(n1830) );
  NOR2X1 U822 ( .A(n1817), .B(n1823), .Y(n1824) );
  NAND2X1 U823 ( .A(n1377), .B(n1376), .Y(n1390) );
  NAND2BX1 U824 ( .AN(n1797), .B(n1796), .Y(n1801) );
  NOR2X1 U825 ( .A(n1788), .B(n1787), .Y(n1797) );
  NOR2X1 U826 ( .A(n1206), .B(n1205), .Y(n1203) );
  NOR2X1 U827 ( .A(n1196), .B(n1199), .Y(n1206) );
  NOR2X1 U828 ( .A(n683), .B(n210), .Y(n1587) );
  AND2X2 U829 ( .A(n1563), .B(n717), .Y(n683) );
  OAI2BB2X1 U830 ( .B0(next_work_cntr[17]), .B1(n2131), .A0N(
        next_work_cntr[17]), .A1N(n2131), .Y(n2142) );
  NAND2BX1 U831 ( .AN(next_work_cntr[16]), .B(n2132), .Y(n2131) );
  NAND2X1 U832 ( .A(n2288), .B(n2287), .Y(n2339) );
  NOR2X1 U833 ( .A(n1764), .B(n1308), .Y(n2288) );
  NOR2X1 U834 ( .A(n1710), .B(n1709), .Y(n1719) );
  OAI31X1 U835 ( .A0(n1711), .A1(n1704), .A2(n1703), .B0(n1702), .Y(n1709) );
  NOR2BX1 U836 ( .AN(n2225), .B(n2224), .Y(n2241) );
  NOR2X1 U837 ( .A(n2216), .B(n2215), .Y(n2224) );
  NOR2X2 U838 ( .A(n827), .B(n830), .Y(n1264) );
  NOR2X1 U839 ( .A(n1755), .B(n2324), .Y(n1763) );
  CLKINVX1 U840 ( .A(n1609), .Y(n1755) );
  NOR2BX1 U841 ( .AN(n1935), .B(n1933), .Y(n1945) );
  NOR2X1 U842 ( .A(n1931), .B(n1930), .Y(n1933) );
  NOR2X1 U843 ( .A(n224), .B(n185), .Y(n882) );
  AND2X4 U844 ( .A(n506), .B(n170), .Y(\DP_OP_665J1_134_4923/I3 ) );
  NOR2BX1 U845 ( .AN(n2280), .B(n2278), .Y(n2315) );
  NOR2X1 U846 ( .A(n1753), .B(n1752), .Y(n1759) );
  NOR2X2 U847 ( .A(n179), .B(n1725), .Y(n1752) );
  NOR2X1 U848 ( .A(n1336), .B(n162), .Y(n1348) );
  NAND2X1 U849 ( .A(N580), .B(N579), .Y(n1336) );
  AOI2BB1X2 U850 ( .A0N(n265), .A1N(n246), .B0(n335), .Y(n594) );
  NAND2X4 U851 ( .A(n664), .B(n170), .Y(n648) );
  NOR2X1 U852 ( .A(n1166), .B(n1170), .Y(n1168) );
  AOI22X1 U853 ( .A0(n1162), .A1(n1161), .B0(n1160), .B1(n1159), .Y(n1170) );
  NOR2X1 U854 ( .A(n2095), .B(n2094), .Y(n2100) );
  OAI21X1 U855 ( .A0(n2093), .A1(n2092), .B0(n2091), .Y(n2094) );
  OAI21X1 U856 ( .A0(n1908), .A1(n1907), .B0(n1906), .Y(n1913) );
  OAI21X1 U857 ( .A0(n1958), .A1(n1805), .B0(n1804), .Y(n1811) );
  NOR2X1 U858 ( .A(n1217), .B(\intadd_3/A[0] ), .Y(n1227) );
  CLKINVX1 U859 ( .A(n1218), .Y(\intadd_3/A[0] ) );
  NOR2X1 U860 ( .A(n1985), .B(n1992), .Y(n1987) );
  OAI21X1 U861 ( .A0(n1980), .A1(n1979), .B0(n1984), .Y(n1992) );
  OAI2BB2X1 U862 ( .B0(n1098), .B1(n1097), .A0N(n1098), .A1N(n1107), .Y(n1114)
         );
  OAI21X1 U863 ( .A0(n1092), .A1(n1088), .B0(n1095), .Y(n1098) );
  NOR2X1 U864 ( .A(n1325), .B(n1327), .Y(n1319) );
  NAND2X2 U865 ( .A(n690), .B(n1306), .Y(n1327) );
  NOR2XL U866 ( .A(n1947), .B(n1899), .Y(n149) );
  CLKINVX1 U867 ( .A(n1896), .Y(n150) );
  OAI21X2 U868 ( .A0(work_cntr[5]), .A1(n946), .B0(n945), .Y(n1947) );
  NOR2XL U869 ( .A(n986), .B(write_addr[18]), .Y(n152) );
  INVXL U870 ( .A(n1055), .Y(n153) );
  AOI211X4 U871 ( .A0(n990), .A1(n151), .B0(n989), .C0(n1354), .Y(n1306) );
  NOR2BX1 U872 ( .AN(n981), .B(n231), .Y(n986) );
  NAND2X1 U873 ( .A(n986), .B(write_addr[18]), .Y(n1055) );
  OAI21X1 U874 ( .A0(n2144), .A1(n2143), .B0(n2145), .Y(n2164) );
  OAI21X1 U875 ( .A0(n2139), .A1(n2138), .B0(n2137), .Y(n2144) );
  OAI21X1 U876 ( .A0(n265), .A1(n162), .B0(n2308), .Y(n638) );
  AOI22X1 U877 ( .A0(n1346), .A1(n718), .B0(n689), .B1(n1345), .Y(n2308) );
  OAI21X1 U878 ( .A0(n1537), .A1(n1540), .B0(n1536), .Y(n1538) );
  OAI21X1 U879 ( .A0(n1019), .A1(n1018), .B0(n1017), .Y(n1032) );
  OAI22X1 U880 ( .A0(n993), .A1(n992), .B0(n1003), .B1(n991), .Y(n1018) );
  NOR2X1 U881 ( .A(curr_time[9]), .B(n413), .Y(n381) );
  NOR2X1 U882 ( .A(n1643), .B(n1633), .Y(n1636) );
  NOR3X1 U883 ( .A(n1632), .B(n1631), .C(n1641), .Y(n1643) );
  NOR4X2 U884 ( .A(n161), .B(n1604), .C(N2666), .D(n1603), .Y(en_photo_num) );
  NOR4X1 U885 ( .A(global_cntr[2]), .B(n1602), .C(n1604), .D(N2666), .Y(n2347)
         );
  CLKINVX1 U886 ( .A(n1515), .Y(n1604) );
  NAND2X1 U887 ( .A(n422), .B(n397), .Y(n420) );
  MXI2X1 U888 ( .A(n438), .B(n396), .S0(curr_time[2]), .Y(n422) );
  NOR3X2 U889 ( .A(n167), .B(n179), .C(n2331), .Y(n1606) );
  NAND2BX1 U890 ( .AN(n1361), .B(n1968), .Y(n1362) );
  CLKINVX1 U891 ( .A(n691), .Y(n1968) );
  OAI21X1 U892 ( .A0(n1283), .A1(n1280), .B0(n1279), .Y(n1298) );
  CLKINVX1 U893 ( .A(n1285), .Y(n1280) );
  OAI2BB2X1 U894 ( .B0(curr_time[12]), .B1(\m_1[3] ), .A0N(curr_time[12]), 
        .A1N(\m_1[3] ), .Y(n936) );
  NAND2X1 U895 ( .A(n315), .B(n319), .Y(\m_1[3] ) );
  NAND2X1 U896 ( .A(n1526), .B(n1580), .Y(n1527) );
  NAND2X1 U897 ( .A(write_cntr[8]), .B(n1580), .Y(n1536) );
  NOR2X1 U898 ( .A(write_cntr[8]), .B(n1580), .Y(n1537) );
  NAND2BX1 U899 ( .AN(n787), .B(n785), .Y(n790) );
  NOR4X2 U900 ( .A(n693), .B(n692), .C(next_glb_cntr[19]), .D(n736), .Y(n2279)
         );
  AOI211X1 U901 ( .A0(n202), .A1(n296), .B0(n297), .C0(n731), .Y(n693) );
  AOI211X1 U902 ( .A0(n201), .A1(n293), .B0(n292), .C0(n731), .Y(n696) );
  NOR2BX2 U903 ( .AN(n726), .B(n729), .Y(n731) );
  NAND2X1 U904 ( .A(n1726), .B(n1728), .Y(n1734) );
  NOR2X1 U905 ( .A(n444), .B(curr_time[17]), .Y(n429) );
  NAND2BX1 U906 ( .AN(n1655), .B(n1656), .Y(n1665) );
  NAND2X1 U907 ( .A(n1646), .B(n1645), .Y(n1656) );
  NOR2X1 U908 ( .A(n307), .B(n306), .Y(n312) );
  NOR2X1 U909 ( .A(write_cntr[6]), .B(n1578), .Y(n1566) );
  NOR2X1 U910 ( .A(N85), .B(n277), .Y(next_work_cntr[0]) );
  NOR2X1 U911 ( .A(n389), .B(n388), .Y(n393) );
  OAI21X1 U912 ( .A0(n1294), .A1(write_addr[10]), .B0(n1241), .Y(n1243) );
  NOR2X1 U913 ( .A(n1295), .B(n244), .Y(n1294) );
  OAI21X1 U914 ( .A0(cr_read_cntr[6]), .A1(n2303), .B0(n973), .Y(n974) );
  OAI22X1 U915 ( .A0(n973), .A1(n2303), .B0(cr_read_cntr[6]), .B1(n972), .Y(
        n975) );
  NOR2X1 U916 ( .A(n249), .B(cr_read_cntr[8]), .Y(n2303) );
  NAND2X1 U917 ( .A(n1306), .B(n1311), .Y(n1322) );
  NOR2X1 U918 ( .A(n164), .B(n1303), .Y(n1311) );
  NOR2X1 U919 ( .A(N2061), .B(n2324), .Y(n1605) );
  CLKINVX1 U920 ( .A(n1374), .Y(n2324) );
  NOR2X1 U921 ( .A(n1347), .B(n2310), .Y(n987) );
  NAND2X1 U922 ( .A(n1348), .B(n272), .Y(n1347) );
  NOR2X1 U923 ( .A(n1388), .B(n1387), .Y(n1382) );
  NOR2X1 U924 ( .A(n2226), .B(n2225), .Y(n2229) );
  OAI211X4 U925 ( .A0(n1614), .A1(n1615), .B0(n1619), .C0(n1613), .Y(n1617) );
  NOR2BX1 U926 ( .AN(n1622), .B(n1618), .Y(n1614) );
  OAI22X2 U927 ( .A0(n776), .A1(n774), .B0(n885), .B1(n208), .Y(n1040) );
  NOR2X1 U928 ( .A(n881), .B(n208), .Y(n776) );
  NOR2X1 U929 ( .A(n2233), .B(n2235), .Y(n2246) );
  OAI21X1 U930 ( .A0(n2232), .A1(n2231), .B0(n2230), .Y(n2235) );
  NOR2X1 U931 ( .A(n161), .B(n1517), .Y(N2664) );
  NAND3X1 U932 ( .A(global_cntr[1]), .B(n1515), .C(n236), .Y(n1517) );
  OAI21X1 U933 ( .A0(curr_time[15]), .A1(n712), .B0(n929), .Y(n931) );
  OAI21X1 U934 ( .A0(curr_time[23]), .A1(n710), .B0(n917), .Y(n919) );
  AOI22X1 U935 ( .A0(n126), .A1(n848), .B0(n125), .B1(n847), .Y(n854) );
  NOR3X1 U936 ( .A(n1148), .B(n1147), .C(n1146), .Y(n1152) );
  OAI2BB2X1 U937 ( .B0(n1130), .B1(n1129), .A0N(n1130), .A1N(n1140), .Y(n1148)
         );
  OAI2BB2X1 U938 ( .B0(n1435), .B1(n1434), .A0N(n1435), .A1N(n1434), .Y(n1440)
         );
  OAI21X1 U939 ( .A0(work_cntr[9]), .A1(n1435), .B0(n1432), .Y(n1437) );
  OAI21X1 U940 ( .A0(n183), .A1(n1431), .B0(n1430), .Y(n1435) );
  OAI21X1 U941 ( .A0(n976), .A1(n977), .B0(cr_read_cntr[4]), .Y(n979) );
  OAI21X1 U942 ( .A0(n975), .A1(n189), .B0(n974), .Y(n977) );
  OAI21X1 U943 ( .A0(n1672), .A1(n214), .B0(n1671), .Y(n1682) );
  OAI22X1 U944 ( .A0(n1015), .A1(n1014), .B0(n1016), .B1(n1013), .Y(n1034) );
  NAND2X2 U945 ( .A(n1017), .B(n1016), .Y(n1231) );
  OAI21X1 U946 ( .A0(n1006), .A1(n1005), .B0(n1004), .Y(n1016) );
  OAI21X1 U947 ( .A0(n176), .A1(n1448), .B0(n1451), .Y(n1456) );
  OAI21X1 U948 ( .A0(n1954), .A1(n1858), .B0(n1862), .Y(n1866) );
  OAI21X1 U949 ( .A0(n1956), .A1(n1876), .B0(n1880), .Y(n1884) );
  OAI31X1 U950 ( .A0(n1822), .A1(n1821), .A2(n1820), .B0(n1819), .Y(n1827) );
  OAI21X1 U951 ( .A0(n1951), .A1(n1810), .B0(n1815), .Y(n1820) );
  OAI211X1 U952 ( .A0(n2337), .A1(n2336), .B0(n2335), .C0(n2334), .Y(
        so_mux_sel[1]) );
  AOI32X4 U953 ( .A0(n776), .A1(n777), .A2(n783), .B0(write_cntr[4]), .B1(n777), .Y(n1771) );
  OAI21X1 U954 ( .A0(n270), .A1(n778), .B0(n885), .Y(n777) );
  OAI22X1 U955 ( .A0(n1562), .A1(n1561), .B0(n1560), .B1(n1559), .Y(n1575) );
  OAI22X1 U956 ( .A0(n1544), .A1(n1543), .B0(n1545), .B1(n1547), .Y(n1560) );
  NAND2X1 U957 ( .A(n1658), .B(n1657), .Y(n1666) );
  OAI22X1 U958 ( .A0(n1653), .A1(n1652), .B0(n1651), .B1(n1650), .Y(n1657) );
  OAI22X1 U959 ( .A0(n1551), .A1(n1550), .B0(n1559), .B1(n1561), .Y(n1577) );
  OAI21X1 U960 ( .A0(n2012), .A1(n2011), .B0(n2010), .Y(n2017) );
  OAI22X1 U961 ( .A0(n2012), .A1(n2004), .B0(n2003), .B1(n2002), .Y(n2013) );
  AOI2BB2X2 U962 ( .B0(n219), .B1(n1988), .A0N(n219), .A1N(n1988), .Y(n2012)
         );
  AOI2BB2X2 U963 ( .B0(n2176), .B1(n2177), .A0N(n2176), .A1N(n2177), .Y(n2197)
         );
  OAI31X4 U964 ( .A0(n2178), .A1(n2172), .A2(n2173), .B0(n2171), .Y(n2177) );
  AOI2BB2X2 U965 ( .B0(n1981), .B1(n2076), .A0N(n1970), .A1N(n181), .Y(n1999)
         );
  NOR2X2 U966 ( .A(work_cntr[15]), .B(n1626), .Y(n1981) );
  OAI31X4 U967 ( .A0(n875), .A1(n1285), .A2(n874), .B0(n873), .Y(n886) );
  NOR2X2 U968 ( .A(n862), .B(n867), .Y(n1285) );
  NAND2BX1 U969 ( .AN(n2248), .B(n2247), .Y(n2256) );
  OAI2BB2X1 U970 ( .B0(n2248), .B1(n2247), .A0N(n2248), .A1N(n2247), .Y(n2254)
         );
  XNOR2X1 U971 ( .A(n423), .B(curr_time[3]), .Y(n418) );
  NAND2X1 U972 ( .A(n394), .B(n393), .Y(n423) );
  MXI2X2 U973 ( .A(n920), .B(curr_time[19]), .S0(n921), .Y(n925) );
  AND2X2 U974 ( .A(n310), .B(n312), .Y(n921) );
  CLKINVX1 U975 ( .A(n1287), .Y(n1301) );
  NOR2X2 U976 ( .A(n876), .B(n886), .Y(n1287) );
  CLKINVX1 U977 ( .A(n1269), .Y(n1268) );
  NAND2X1 U978 ( .A(n848), .B(n1269), .Y(n847) );
  OAI22X1 U979 ( .A0(n1272), .A1(n1271), .B0(n1270), .B1(n1269), .Y(n1275) );
  AOI32X1 U980 ( .A0(N85), .A1(n688), .A2(n2327), .B0(n2337), .B1(n688), .Y(
        n2336) );
  NAND2X1 U981 ( .A(n688), .B(curr_photo_size[1]), .Y(n2330) );
  AND2X2 U982 ( .A(n329), .B(n328), .Y(n688) );
  MXI2X2 U983 ( .A(n377), .B(n937), .S0(n379), .Y(n411) );
  OAI21X1 U984 ( .A0(n935), .A1(n936), .B0(n372), .Y(n379) );
  NAND2BX1 U985 ( .AN(n1681), .B(n1680), .Y(n1697) );
  OAI2BB2X1 U986 ( .B0(next_work_cntr[14]), .B1(n2128), .A0N(
        next_work_cntr[14]), .A1N(n2128), .Y(n2151) );
  NOR2X1 U987 ( .A(n2128), .B(next_work_cntr[14]), .Y(n2140) );
  OAI2BB2X2 U988 ( .B0(n219), .B1(n953), .A0N(n219), .A1N(n953), .Y(n1951) );
  NOR2X1 U989 ( .A(next_work_cntr[7]), .B(n2203), .Y(n2191) );
  OAI2BB2X1 U990 ( .B0(next_work_cntr[7]), .B1(n2203), .A0N(next_work_cntr[7]), 
        .A1N(n2203), .Y(n2216) );
  CLKINVX1 U991 ( .A(n1877), .Y(n1956) );
  CLKINVX1 U992 ( .A(n1248), .Y(n1249) );
  NOR2X1 U993 ( .A(n1248), .B(n792), .Y(n794) );
  OAI2BB2X1 U994 ( .B0(n1569), .B1(n1568), .A0N(n1569), .A1N(n1568), .Y(n1597)
         );
  NOR2X2 U995 ( .A(n1554), .B(n1552), .Y(n1569) );
  NOR2X1 U996 ( .A(write_cntr[7]), .B(n1579), .Y(n1552) );
  CLKINVX1 U997 ( .A(n1540), .Y(n1554) );
  NAND2BX1 U998 ( .AN(next_work_cntr[6]), .B(n2217), .Y(n2203) );
  NOR2X1 U999 ( .A(n277), .B(n1948), .Y(next_work_cntr[6]) );
  NOR2BX1 U1000 ( .AN(n2140), .B(next_work_cntr[15]), .Y(n2132) );
  CLKINVX1 U1001 ( .A(n1798), .Y(n1958) );
  NOR2X1 U1002 ( .A(next_work_cntr[9]), .B(n2123), .Y(n2124) );
  CLKINVX1 U1003 ( .A(n1859), .Y(n1954) );
  NAND2X1 U1004 ( .A(n154), .B(n155), .Y(n1571) );
  CLKINVX1 U1005 ( .A(n1555), .Y(n156) );
  INVXL U1006 ( .A(n1556), .Y(n157) );
  NAND2XL U1007 ( .A(n1556), .B(n1555), .Y(n154) );
  NAND2X1 U1008 ( .A(n156), .B(n157), .Y(n155) );
  OAI21X1 U1009 ( .A0(n1554), .A1(n1565), .B0(n1553), .Y(n1555) );
  OAI2BB2X1 U1010 ( .B0(n1571), .B1(n1570), .A0N(n1571), .A1N(n1570), .Y(n1596) );
  NOR2BX2 U1011 ( .AN(n1536), .B(n1537), .Y(n1556) );
  AOI2BB2X2 U1012 ( .B0(n1539), .B1(n1538), .A0N(n1539), .A1N(n1538), .Y(n1558) );
  NAND3X1 U1013 ( .A(write_cntr[8]), .B(write_cntr[10]), .C(n1539), .Y(n1526)
         );
  NOR2BX2 U1014 ( .AN(n1523), .B(n1524), .Y(n1539) );
  NOR2BX2 U1015 ( .AN(n2163), .B(n2158), .Y(n2169) );
  OAI21X1 U1016 ( .A0(n2156), .A1(n2152), .B0(n2151), .Y(n2163) );
  OAI21X2 U1017 ( .A0(work_cntr[8]), .A1(n947), .B0(n948), .Y(n1949) );
  NAND2X1 U1018 ( .A(work_cntr[8]), .B(n947), .Y(n948) );
  NOR2X1 U1019 ( .A(n176), .B(n944), .Y(n947) );
  AOI2BB2X2 U1020 ( .B0(n2159), .B1(n2160), .A0N(n2159), .A1N(n2160), .Y(n2175) );
  NOR2BX1 U1021 ( .AN(n2160), .B(n2159), .Y(n2168) );
  OAI2BB2X2 U1022 ( .B0(n2127), .B1(n2126), .A0N(n2127), .A1N(n2126), .Y(n2159) );
  AOI32X4 U1023 ( .A0(n2136), .A1(n2148), .A2(n2135), .B0(n2134), .B1(n2148), 
        .Y(n2155) );
  OAI211X4 U1024 ( .A0(n2133), .A1(n2136), .B0(n2141), .C0(n2134), .Y(n2148)
         );
  CLKINVX1 U1025 ( .A(n1775), .Y(n1027) );
  AOI32X4 U1026 ( .A0(n210), .A1(n783), .A2(n778), .B0(n777), .B1(
        write_cntr[5]), .Y(n1775) );
  NAND2X1 U1027 ( .A(n982), .B(write_addr[11]), .Y(n983) );
  OAI21X1 U1028 ( .A0(n982), .A1(write_addr[11]), .B0(n983), .Y(n1292) );
  NAND2X1 U1029 ( .A(write_addr[11]), .B(n1289), .Y(n1303) );
  CLKINVX1 U1030 ( .A(n1934), .Y(n1939) );
  AOI21X1 U1031 ( .A0(write_cntr[4]), .A1(n1767), .B0(n1587), .Y(n1593) );
  AND2X2 U1032 ( .A(n1767), .B(n383), .Y(n458) );
  NOR2X2 U1033 ( .A(n1767), .B(n404), .Y(n464) );
  NAND2X2 U1034 ( .A(n362), .B(n1583), .Y(n1767) );
  AND2X2 U1035 ( .A(n911), .B(n907), .Y(n1240) );
  OAI21X1 U1036 ( .A0(cr_read_cntr[6]), .A1(n2299), .B0(n2298), .Y(n2301) );
  CLKINVX1 U1037 ( .A(n2299), .Y(n2302) );
  NOR2BX1 U1038 ( .AN(n2293), .B(n2299), .Y(n2294) );
  NAND2X2 U1039 ( .A(n2289), .B(next_en_si), .Y(n2299) );
  NOR3X2 U1040 ( .A(work_cntr[17]), .B(work_cntr[18]), .C(n1982), .Y(n1975) );
  CLKINVX1 U1041 ( .A(n1975), .Y(n1971) );
  AOI22X1 U1042 ( .A0(n1976), .A1(work_cntr[18]), .B0(n1975), .B1(n2076), .Y(
        n1979) );
  OAI21X2 U1043 ( .A0(n1975), .A1(n212), .B0(n1755), .Y(n1615) );
  NAND2X1 U1044 ( .A(write_cntr[13]), .B(write_cntr[12]), .Y(n751) );
  NAND2X1 U1045 ( .A(write_addr[15]), .B(write_addr[14]), .Y(n1358) );
  OAI22X1 U1046 ( .A0(write_addr[14]), .A1(n1314), .B0(n246), .B1(n1310), .Y(
        n1312) );
  OAI22X1 U1047 ( .A0(n1770), .A1(n1288), .B0(n898), .B1(\intadd_4/A[1] ), .Y(
        n909) );
  NOR2X2 U1048 ( .A(n893), .B(n897), .Y(n1288) );
  NOR2X2 U1049 ( .A(n1967), .B(n277), .Y(next_work_cntr[19]) );
  CLKINVX1 U1050 ( .A(n641), .Y(n655) );
  NAND2X4 U1051 ( .A(n664), .B(read_cntr[0]), .Y(n641) );
  NOR2X2 U1052 ( .A(n1601), .B(n371), .Y(n463) );
  NOR2X1 U1053 ( .A(n277), .B(n1950), .Y(next_work_cntr[16]) );
  OA21X1 U1054 ( .A0(n1950), .A1(n1796), .B0(n1790), .Y(n1800) );
  OAI21X1 U1055 ( .A0(n1797), .A1(n1789), .B0(n1950), .Y(n1790) );
  OAI21X2 U1056 ( .A0(work_cntr[16]), .A1(n955), .B0(n1783), .Y(n1950) );
  NAND2X1 U1057 ( .A(work_cntr[16]), .B(n955), .Y(n1783) );
  NOR3X2 U1058 ( .A(n181), .B(n219), .C(n953), .Y(n955) );
  OAI21X2 U1059 ( .A0(n885), .A1(n203), .B0(n760), .Y(n961) );
  OAI21X2 U1060 ( .A0(n984), .A1(write_addr[13]), .B0(n1310), .Y(n1323) );
  NAND2X1 U1061 ( .A(n984), .B(write_addr[13]), .Y(n1310) );
  NOR2X1 U1062 ( .A(n983), .B(n164), .Y(n984) );
  NAND2BX1 U1063 ( .AN(n1323), .B(n1311), .Y(n1317) );
  NOR3X1 U1064 ( .A(n1358), .B(n1323), .C(n1322), .Y(n1324) );
  NOR2X2 U1065 ( .A(n277), .B(n1955), .Y(next_work_cntr[11]) );
  OAI21X1 U1066 ( .A0(n1955), .A1(n1845), .B0(n1844), .Y(n1850) );
  OAI21X2 U1067 ( .A0(work_cntr[11]), .A1(n950), .B0(n951), .Y(n1955) );
  NAND2X1 U1068 ( .A(work_cntr[11]), .B(n950), .Y(n951) );
  NOR3X2 U1069 ( .A(n183), .B(n214), .C(n948), .Y(n950) );
  NOR3BX1 U1070 ( .AN(n2176), .B(n2175), .C(n2186), .Y(n2178) );
  NOR3X1 U1071 ( .A(n2183), .B(n2197), .C(n2186), .Y(n2187) );
  OAI21X2 U1072 ( .A0(n2167), .A1(n2166), .B0(n2170), .Y(n2186) );
  NOR3X1 U1073 ( .A(n1710), .B(n1707), .C(n1717), .Y(n1711) );
  OAI21X2 U1074 ( .A0(n1686), .A1(n1685), .B0(n1690), .Y(n1707) );
  NAND2X2 U1075 ( .A(n1164), .B(n2119), .Y(n1911) );
  CLKINVX1 U1076 ( .A(n1606), .Y(n2119) );
  CLKINVX1 U1077 ( .A(n1274), .Y(n1277) );
  NOR2X2 U1078 ( .A(n850), .B(n854), .Y(n1274) );
  OAI22X2 U1079 ( .A0(work_cntr[4]), .A1(n1164), .B0(n180), .B1(n1163), .Y(
        n1177) );
  CLKINVX1 U1080 ( .A(n1163), .Y(n1164) );
  NOR2X2 U1081 ( .A(N2063), .B(n957), .Y(n1163) );
  INVX3 U1082 ( .A(n1776), .Y(n1023) );
  OAI221X4 U1083 ( .A0(n783), .A1(write_cntr[6]), .B0(n780), .B1(write_cntr[6]), .C0(n781), .Y(n1776) );
  OAI21X1 U1084 ( .A0(n2120), .A1(n1929), .B0(n1928), .Y(n1938) );
  AOI21X2 U1085 ( .A0(n2331), .A1(N2062), .B0(n2322), .Y(n2120) );
  NOR2X1 U1086 ( .A(n2331), .B(N2062), .Y(n2322) );
  INVX3 U1087 ( .A(n773), .Y(n885) );
  OAI21X2 U1088 ( .A0(n1056), .A1(write_addr[8]), .B0(n1295), .Y(n1297) );
  NAND2X1 U1089 ( .A(n1056), .B(write_addr[8]), .Y(n1295) );
  CLKINVX1 U1090 ( .A(n1356), .Y(n1056) );
  NOR2X1 U1091 ( .A(n244), .B(n1297), .Y(n1296) );
  NOR2X2 U1092 ( .A(work_cntr[5]), .B(work_cntr[4]), .Y(n2057) );
  OAI22X1 U1093 ( .A0(n1257), .A1(n826), .B0(n825), .B1(n824), .Y(n830) );
  CLKINVX1 U1094 ( .A(n1257), .Y(n1256) );
  NOR2X1 U1095 ( .A(n1257), .B(n1259), .Y(n1261) );
  NOR2X2 U1096 ( .A(n815), .B(n816), .Y(n1257) );
  AOI32X4 U1097 ( .A0(n1777), .A1(n783), .A2(n782), .B0(n781), .B1(
        write_cntr[7]), .Y(n1778) );
  CLKINVX2 U1098 ( .A(n270), .Y(n783) );
  AOI22X2 U1099 ( .A0(n1053), .A1(n1052), .B0(n1051), .B1(n1050), .Y(
        \intadd_3/B[0] ) );
  CLKINVX1 U1100 ( .A(next_cr_x[6]), .Y(n1230) );
  INVX3 U1101 ( .A(n770), .Y(next_cr_x[6]) );
  AOI222X4 U1102 ( .A0(n967), .A1(n1223), .B0(n967), .B1(n966), .C0(n965), 
        .C1(next_cr_x[5]), .Y(n993) );
  NAND2X2 U1103 ( .A(n969), .B(n968), .Y(next_cr_x[5]) );
  CLKINVX1 U1104 ( .A(n1355), .Y(n718) );
  NAND2X2 U1105 ( .A(n1330), .B(n690), .Y(n1355) );
  INVX3 U1106 ( .A(n645), .Y(n647) );
  NAND2X2 U1107 ( .A(n158), .B(n159), .Y(n964) );
  CLKINVX1 U1108 ( .A(n758), .Y(n160) );
  NAND2XL U1109 ( .A(n160), .B(n107), .Y(n158) );
  NAND2X1 U1110 ( .A(n160), .B(n885), .Y(n159) );
  AOI2BB2X2 U1111 ( .B0(n964), .B1(n963), .A0N(n964), .A1N(n963), .Y(n1001) );
  NOR3X1 U1112 ( .A(n115), .B(n998), .C(n964), .Y(n966) );
  NOR2X1 U1113 ( .A(n1779), .B(n964), .Y(n768) );
  INVX3 U1114 ( .A(n1372), .Y(n571) );
  OAI211X4 U1115 ( .A0(n1369), .A1(n1368), .B0(n1367), .C0(n1366), .Y(n1372)
         );
  CLKBUFX8 U1116 ( .A(n686), .Y(n273) );
  CLKINVX1 U1117 ( .A(n2314), .Y(n686) );
  NAND2X4 U1118 ( .A(n1368), .B(n657), .Y(n649) );
  CLKINVX1 U1119 ( .A(n2077), .Y(n2076) );
  NAND2X4 U1120 ( .A(n179), .B(n2097), .Y(n2077) );
  AND2X4 U1121 ( .A(read_cntr[0]), .B(n506), .Y(\DP_OP_665J1_134_4923/I4 ) );
  NOR2X1 U1122 ( .A(n685), .B(n505), .Y(n506) );
  INVX4 U1123 ( .A(n169), .Y(n269) );
  NOR2X6 U1124 ( .A(n266), .B(n573), .Y(\DP_OP_665J1_134_4923/I7 ) );
  BUFX4 U1125 ( .A(n662), .Y(n266) );
  INVX6 U1126 ( .A(n171), .Y(n276) );
  NOR3X6 U1127 ( .A(n504), .B(n685), .C(n572), .Y(\DP_OP_665J1_134_4923/I2 )
         );
  AND2X2 U1128 ( .A(\next_write_addr_w[0] ), .B(n1056), .Y(n685) );
  INVXL U1129 ( .A(n279), .Y(n1603) );
  NOR2X1 U1130 ( .A(global_cntr[1]), .B(global_cntr[0]), .Y(n279) );
  NOR2X2 U1131 ( .A(global_cntr[2]), .B(n1517), .Y(N2622) );
  NAND3X2 U1132 ( .A(n28), .B(n172), .C(n205), .Y(N2666) );
  XOR2XL U1133 ( .A(curr_photo[0]), .B(curr_photo[1]), .Y(n366) );
  NAND2XL U1134 ( .A(n2316), .B(n2315), .Y(n2320) );
  INVXL U1135 ( .A(n2192), .Y(next_work_cntr[8]) );
  NOR2XL U1136 ( .A(n2120), .B(n277), .Y(next_work_cntr[2]) );
  NOR2XL U1137 ( .A(n277), .B(n1908), .Y(next_work_cntr[4]) );
  NOR2XL U1138 ( .A(n1911), .B(n277), .Y(next_work_cntr[3]) );
  NOR2BXL U1139 ( .AN(N1235), .B(n2334), .Y(n2346) );
  NOR2BXL U1140 ( .AN(N1236), .B(n2334), .Y(n2345) );
  NOR2BXL U1141 ( .AN(N1237), .B(n2334), .Y(n2344) );
  NOR2BXL U1142 ( .AN(N1238), .B(n2334), .Y(n2343) );
  NOR2BXL U1143 ( .AN(N1239), .B(n2334), .Y(n2342) );
  NAND2XL U1144 ( .A(n464), .B(n432), .Y(n433) );
  NAND2BXL U1145 ( .AN(n928), .B(n429), .Y(n430) );
  INVXL U1146 ( .A(n429), .Y(n431) );
  AOI211XL U1147 ( .A0(n428), .A1(n427), .B0(n426), .C0(n425), .Y(n434) );
  NOR2XL U1148 ( .A(n921), .B(n417), .Y(n426) );
  INVXL U1149 ( .A(n463), .Y(n417) );
  INVXL U1150 ( .A(n381), .Y(n415) );
  INVXL U1151 ( .A(n411), .Y(n416) );
  INVXL U1152 ( .A(n465), .Y(n428) );
  OAI211XL U1153 ( .A0(curr_time[17]), .A1(n446), .B0(n464), .C0(n445), .Y(
        n447) );
  NAND2XL U1154 ( .A(curr_time[17]), .B(n454), .Y(n445) );
  INVXL U1155 ( .A(n444), .Y(n446) );
  AOI211XL U1156 ( .A0(n463), .A1(h_1[1]), .B0(n443), .C0(n442), .Y(n448) );
  INVXL U1157 ( .A(n438), .Y(n439) );
  AOI21XL U1158 ( .A0(n451), .A1(curr_time[1]), .B0(n437), .Y(n441) );
  NOR2XL U1159 ( .A(n436), .B(n465), .Y(n443) );
  XOR2XL U1160 ( .A(n457), .B(curr_time[9]), .Y(n436) );
  INVXL U1161 ( .A(n435), .Y(n449) );
  INVXL U1162 ( .A(n450), .Y(n461) );
  NAND2XL U1163 ( .A(n464), .B(\h_0[0] ), .Y(n455) );
  AOI211XL U1164 ( .A0(n463), .A1(n454), .B0(n453), .C0(n452), .Y(n456) );
  NOR2XL U1165 ( .A(n683), .B(n1768), .Y(n383) );
  INVXL U1166 ( .A(n399), .Y(n402) );
  INVXL U1167 ( .A(curr_time[1]), .Y(n397) );
  NOR2XL U1168 ( .A(n400), .B(n401), .Y(n396) );
  INVXL U1169 ( .A(n395), .Y(n401) );
  NAND2XL U1170 ( .A(n418), .B(n398), .Y(n399) );
  NOR2XL U1171 ( .A(n393), .B(n942), .Y(n390) );
  AOI21XL U1172 ( .A0(n423), .A1(n715), .B0(n943), .Y(n391) );
  INVXL U1173 ( .A(n387), .Y(n388) );
  NOR2XL U1174 ( .A(n386), .B(n385), .Y(n389) );
  INVXL U1175 ( .A(curr_time[6]), .Y(n385) );
  NAND2XL U1176 ( .A(n943), .B(n715), .Y(n942) );
  INVXL U1177 ( .A(curr_time[3]), .Y(n715) );
  NOR2XL U1178 ( .A(curr_time[5]), .B(curr_time[6]), .Y(n940) );
  NAND3XL U1179 ( .A(n386), .B(curr_time[6]), .C(n322), .Y(n323) );
  NAND2BXL U1180 ( .AN(curr_time[5]), .B(curr_time[7]), .Y(n322) );
  NAND2BXL U1181 ( .AN(n941), .B(n384), .Y(n386) );
  INVXL U1182 ( .A(curr_time[4]), .Y(n384) );
  NAND3XL U1183 ( .A(curr_time[7]), .B(curr_time[6]), .C(n714), .Y(n939) );
  INVXL U1184 ( .A(curr_time[5]), .Y(n714) );
  INVXL U1185 ( .A(curr_time[2]), .Y(n398) );
  NOR2BXL U1186 ( .AN(\m_0[0] ), .B(n465), .Y(n453) );
  INVXL U1187 ( .A(n927), .Y(n405) );
  NAND2XL U1188 ( .A(n410), .B(n313), .Y(n927) );
  NAND2XL U1189 ( .A(n406), .B(n410), .Y(h_1[1]) );
  NAND2XL U1190 ( .A(n925), .B(n711), .Y(n926) );
  NOR2XL U1191 ( .A(curr_time[19]), .B(n921), .Y(n923) );
  INVXL U1192 ( .A(n922), .Y(n308) );
  NAND2XL U1193 ( .A(n924), .B(n920), .Y(n922) );
  INVXL U1194 ( .A(curr_time[19]), .Y(n920) );
  NAND3XL U1195 ( .A(n304), .B(curr_time[22]), .C(n300), .Y(n301) );
  NAND2BXL U1196 ( .AN(curr_time[21]), .B(curr_time[23]), .Y(n300) );
  INVXL U1197 ( .A(n312), .Y(n309) );
  INVXL U1198 ( .A(n305), .Y(n306) );
  NOR2XL U1199 ( .A(n304), .B(n303), .Y(n307) );
  INVXL U1200 ( .A(curr_time[22]), .Y(n303) );
  NAND2BXL U1201 ( .AN(n919), .B(n302), .Y(n304) );
  INVXL U1202 ( .A(curr_time[20]), .Y(n302) );
  NAND3XL U1203 ( .A(curr_time[23]), .B(curr_time[22]), .C(n710), .Y(n917) );
  INVXL U1204 ( .A(curr_time[21]), .Y(n710) );
  INVXL U1205 ( .A(curr_time[17]), .Y(n408) );
  INVXL U1206 ( .A(n459), .Y(n371) );
  NAND3XL U1207 ( .A(n403), .B(n683), .C(n370), .Y(n404) );
  INVXL U1208 ( .A(n1768), .Y(n370) );
  NOR3XL U1209 ( .A(n1580), .B(n1579), .C(n1578), .Y(n1581) );
  OAI211XL U1210 ( .A0(n1598), .A1(n1597), .B0(n1596), .C0(n1595), .Y(n1599)
         );
  INVXL U1211 ( .A(n1588), .Y(n1591) );
  INVXL U1212 ( .A(n1585), .Y(n1574) );
  INVXL U1213 ( .A(n1584), .Y(n362) );
  NAND2XL U1214 ( .A(n1586), .B(n1585), .Y(n1598) );
  NOR2XL U1215 ( .A(n1571), .B(n1570), .Y(n1572) );
  NAND2XL U1216 ( .A(n1577), .B(n1576), .Y(n1563) );
  NOR2XL U1217 ( .A(n1558), .B(n1557), .Y(n1550) );
  NAND3XL U1218 ( .A(write_cntr[5]), .B(n1569), .C(n1588), .Y(n1564) );
  INVXL U1219 ( .A(n1552), .Y(n1553) );
  INVXL U1220 ( .A(n1575), .Y(n717) );
  INVXL U1221 ( .A(n1546), .Y(n1548) );
  NAND2XL U1222 ( .A(write_cntr[7]), .B(n1579), .Y(n1540) );
  INVXL U1223 ( .A(n1560), .Y(n1562) );
  NOR2XL U1224 ( .A(n1542), .B(n1541), .Y(n1543) );
  INVXL U1225 ( .A(n1532), .Y(n1534) );
  NOR2XL U1226 ( .A(n130), .B(n1527), .Y(n1529) );
  NAND3XL U1227 ( .A(write_cntr[7]), .B(n1539), .C(n1556), .Y(n1535) );
  OAI2BB2XL U1228 ( .B0(write_cntr[11]), .B1(n1520), .A0N(write_cntr[11]), 
        .A1N(n1520), .Y(n1528) );
  NAND2XL U1229 ( .A(write_cntr[10]), .B(n260), .Y(n1520) );
  INVXL U1230 ( .A(n1523), .Y(n260) );
  INVXL U1231 ( .A(n938), .Y(n376) );
  NAND2XL U1232 ( .A(n435), .B(n713), .Y(n378) );
  NOR2XL U1233 ( .A(curr_time[11]), .B(n933), .Y(n935) );
  INVXL U1234 ( .A(n377), .Y(n380) );
  NAND2XL U1235 ( .A(n936), .B(n932), .Y(n934) );
  INVXL U1236 ( .A(curr_time[11]), .Y(n932) );
  NAND3XL U1237 ( .A(n318), .B(curr_time[14]), .C(n314), .Y(n315) );
  NAND2BXL U1238 ( .AN(curr_time[13]), .B(curr_time[15]), .Y(n314) );
  INVXL U1239 ( .A(n319), .Y(n320) );
  NOR2XL U1240 ( .A(curr_time[13]), .B(curr_time[14]), .Y(n930) );
  NOR2XL U1241 ( .A(n318), .B(n317), .Y(n321) );
  INVXL U1242 ( .A(curr_time[14]), .Y(n317) );
  NAND2BXL U1243 ( .AN(n931), .B(n316), .Y(n318) );
  INVXL U1244 ( .A(curr_time[12]), .Y(n316) );
  NAND3XL U1245 ( .A(curr_time[15]), .B(curr_time[14]), .C(n712), .Y(n929) );
  INVXL U1246 ( .A(curr_time[13]), .Y(n712) );
  NAND2XL U1247 ( .A(n979), .B(n980), .Y(n470) );
  MXI2XL U1248 ( .A(cr_read_cntr[4]), .B(n979), .S0(n980), .Y(n502) );
  AND2XL U1249 ( .A(n500), .B(cr_read_cntr[3]), .Y(n503) );
  NAND2XL U1250 ( .A(n979), .B(n469), .Y(n500) );
  INVXL U1251 ( .A(n978), .Y(n468) );
  AND2XL U1252 ( .A(n975), .B(n189), .Y(n976) );
  NAND2XL U1253 ( .A(n972), .B(cr_read_cntr[6]), .Y(n973) );
  NAND2XL U1254 ( .A(n249), .B(cr_read_cntr[8]), .Y(n972) );
  MXI2XL U1255 ( .A(n2339), .B(n2338), .S0(read_cntr[0]), .Y(n519) );
  NAND2XL U1256 ( .A(n2340), .B(n2339), .Y(n2338) );
  INVXL U1257 ( .A(n658), .Y(n360) );
  OAI211XL U1258 ( .A0(n1760), .A1(n1748), .B0(n1747), .C0(n1746), .Y(n1749)
         );
  NAND2XL U1259 ( .A(n1760), .B(n1748), .Y(n1746) );
  NAND2XL U1260 ( .A(n1745), .B(n1744), .Y(n1748) );
  NOR2BXL U1261 ( .AN(n2323), .B(n1751), .Y(n1740) );
  NAND2XL U1262 ( .A(n681), .B(n2328), .Y(n2329) );
  NAND2BXL U1263 ( .AN(n2326), .B(n2325), .Y(n2337) );
  INVXL U1264 ( .A(n2321), .Y(n2325) );
  NAND2XL U1265 ( .A(n273), .B(write_addr[15]), .Y(n333) );
  NAND2XL U1266 ( .A(n273), .B(n271), .Y(n357) );
  NAND2XL U1267 ( .A(write_addr[14]), .B(n273), .Y(n336) );
  NAND2XL U1268 ( .A(n273), .B(write_addr[16]), .Y(n356) );
  MXI2XL U1269 ( .A(n2299), .B(n682), .S0(N1232), .Y(n499) );
  AOI211XL U1270 ( .A0(n2292), .A1(n257), .B0(n2299), .C0(n2293), .Y(n364) );
  NAND2XL U1271 ( .A(n273), .B(\next_write_addr_w[0] ), .Y(n359) );
  AOI21XL U1272 ( .A0(n249), .A1(n2304), .B0(n2306), .Y(n492) );
  NAND2XL U1273 ( .A(cr_read_cntr[6]), .B(n2300), .Y(n2304) );
  INVXL U1274 ( .A(n2303), .Y(n2305) );
  NAND2XL U1275 ( .A(cr_read_cntr[5]), .B(cr_read_cntr[4]), .Y(n2297) );
  OAI211XL U1276 ( .A0(n2282), .A1(next_glb_cntr[2]), .B0(n2281), .C0(n2280), 
        .Y(n2283) );
  OAI21X1 U1277 ( .A0(global_cntr[2]), .A1(n1602), .B0(n1516), .Y(
        next_glb_cntr[2]) );
  INVXL U1278 ( .A(n2279), .Y(n2282) );
  OAI211XL U1279 ( .A0(n2273), .A1(n2272), .B0(n2271), .C0(n2270), .Y(n2274)
         );
  MXI2XL U1280 ( .A(n2273), .B(n2272), .S0(n2269), .Y(n2270) );
  NOR2XL U1281 ( .A(N2061), .B(n277), .Y(n2269) );
  NOR2XL U1282 ( .A(n2268), .B(n2267), .Y(n2271) );
  NAND2XL U1283 ( .A(si_sel), .B(next_work_cntr[0]), .Y(n2267) );
  INVXL U1284 ( .A(n2266), .Y(n2272) );
  NAND2XL U1285 ( .A(n2262), .B(n2261), .Y(n2258) );
  NAND2XL U1286 ( .A(n2257), .B(n2256), .Y(n2255) );
  INVXL U1287 ( .A(n2260), .Y(n2253) );
  NAND2XL U1288 ( .A(n2250), .B(n2249), .Y(n2264) );
  INVXL U1289 ( .A(n2254), .Y(n2265) );
  INVXL U1290 ( .A(n2252), .Y(n2249) );
  INVXL U1291 ( .A(n2237), .Y(n2239) );
  INVXL U1292 ( .A(n2234), .Y(n2238) );
  INVXL U1293 ( .A(n2227), .Y(n2228) );
  NAND2XL U1294 ( .A(n2226), .B(n2225), .Y(n2231) );
  AOI211XL U1295 ( .A0(n2233), .A1(n2237), .B0(n2224), .C0(n2234), .Y(n2232)
         );
  NOR2XL U1296 ( .A(n2226), .B(n2227), .Y(n2221) );
  NAND2XL U1297 ( .A(n2241), .B(n2223), .Y(n2227) );
  OAI211XL U1298 ( .A0(n2216), .A1(n2220), .B0(n2210), .C0(n2209), .Y(n2211)
         );
  INVXL U1299 ( .A(n2206), .Y(n2207) );
  INVXL U1300 ( .A(n2212), .Y(n2214) );
  NAND2BXL U1301 ( .AN(n2205), .B(n2204), .Y(n2212) );
  NAND2XL U1302 ( .A(n2194), .B(n2193), .Y(n2210) );
  INVXL U1303 ( .A(n2187), .Y(n2188) );
  NOR2BXL U1304 ( .AN(n2196), .B(n2197), .Y(n2190) );
  INVXL U1305 ( .A(n2178), .Y(n2179) );
  NOR2XL U1306 ( .A(n2185), .B(n2186), .Y(n2180) );
  AOI21XL U1307 ( .A0(n2175), .A1(n2174), .B0(n2173), .Y(n2181) );
  NAND2XL U1308 ( .A(n2166), .B(n2167), .Y(n2174) );
  NAND2XL U1309 ( .A(n2169), .B(n2168), .Y(n2162) );
  AOI21XL U1310 ( .A0(n2155), .A1(n2154), .B0(n2153), .Y(n2157) );
  AOI21XL U1311 ( .A0(n2148), .A1(n2147), .B0(n2146), .Y(n2150) );
  NAND2XL U1312 ( .A(n2142), .B(n2141), .Y(n2147) );
  NAND2XL U1313 ( .A(n2144), .B(n2143), .Y(n2154) );
  NAND3XL U1314 ( .A(n2139), .B(n2141), .C(n2138), .Y(n2137) );
  INVXL U1315 ( .A(n2146), .Y(n2139) );
  INVXL U1316 ( .A(n2135), .Y(n2133) );
  NAND2XL U1317 ( .A(n2138), .B(n2142), .Y(n2135) );
  INVXL U1318 ( .A(n2183), .Y(n2182) );
  INVXL U1319 ( .A(n2236), .Y(n2233) );
  NAND4XL U1320 ( .A(n2268), .B(si_sel), .C(next_work_cntr[0]), .D(n2121), .Y(
        n2276) );
  XOR2XL U1321 ( .A(n2109), .B(n2108), .Y(n2110) );
  INVXL U1322 ( .A(n2094), .Y(n2103) );
  AND3XL U1323 ( .A(n2095), .B(n2091), .C(n2102), .Y(n2098) );
  NAND3XL U1324 ( .A(n2093), .B(n2092), .C(n2090), .Y(n2091) );
  INVXL U1325 ( .A(n2089), .Y(n2093) );
  INVXL U1326 ( .A(n2083), .Y(n2085) );
  NAND3XL U1327 ( .A(n2075), .B(n2082), .C(n2078), .Y(n2090) );
  NAND3XL U1328 ( .A(n2080), .B(n2079), .C(n2074), .Y(n2078) );
  INVXL U1329 ( .A(n2073), .Y(n2080) );
  INVXL U1330 ( .A(n2081), .Y(n2075) );
  INVXL U1331 ( .A(n2067), .Y(n2069) );
  NOR2XL U1332 ( .A(work_cntr[4]), .B(n2077), .Y(n2061) );
  NOR2XL U1333 ( .A(n2060), .B(n2077), .Y(n2059) );
  INVXL U1334 ( .A(n2057), .Y(n2060) );
  INVXL U1335 ( .A(n2071), .Y(n2072) );
  NAND3XL U1336 ( .A(n2056), .B(n2066), .C(n2062), .Y(n2074) );
  NAND3XL U1337 ( .A(n2064), .B(n2063), .C(n2055), .Y(n2062) );
  INVXL U1338 ( .A(n2054), .Y(n2064) );
  INVXL U1339 ( .A(n2065), .Y(n2056) );
  INVXL U1340 ( .A(n2048), .Y(n2050) );
  NOR2XL U1341 ( .A(n2058), .B(n2077), .Y(n2042) );
  INVXL U1342 ( .A(n2052), .Y(n2053) );
  NAND3XL U1343 ( .A(n2039), .B(n2047), .C(n2043), .Y(n2055) );
  NAND3XL U1344 ( .A(n2045), .B(n2044), .C(n2038), .Y(n2043) );
  INVXL U1345 ( .A(n2037), .Y(n2045) );
  INVXL U1346 ( .A(n2046), .Y(n2039) );
  INVXL U1347 ( .A(n2031), .Y(n2033) );
  INVXL U1348 ( .A(n2035), .Y(n2036) );
  NAND3XL U1349 ( .A(n2023), .B(n2030), .C(n2026), .Y(n2038) );
  NAND3XL U1350 ( .A(n2028), .B(n2027), .C(n2022), .Y(n2026) );
  INVXL U1351 ( .A(n2029), .Y(n2023) );
  INVXL U1352 ( .A(n2017), .Y(n2015) );
  INVXL U1353 ( .A(n2019), .Y(n2020) );
  INVXL U1354 ( .A(n2013), .Y(n2006) );
  NAND2XL U1355 ( .A(n1997), .B(n1996), .Y(n2001) );
  INVXL U1356 ( .A(n1992), .Y(n1995) );
  NAND2XL U1357 ( .A(n1991), .B(n1990), .Y(n1997) );
  NOR2XL U1358 ( .A(work_cntr[12]), .B(n2007), .Y(n1989) );
  NOR2XL U1359 ( .A(n2009), .B(n2003), .Y(n2004) );
  AND2XL U1360 ( .A(n1998), .B(n1999), .Y(n2003) );
  INVXL U1361 ( .A(n1993), .Y(n1990) );
  NOR2BXL U1362 ( .AN(n1981), .B(n2077), .Y(n1983) );
  AND2XL U1363 ( .A(n1980), .B(n1979), .Y(n1985) );
  NAND2XL U1364 ( .A(n2076), .B(n1973), .Y(n1976) );
  NOR2XL U1365 ( .A(n1982), .B(n2077), .Y(n1974) );
  NOR2XL U1366 ( .A(n1971), .B(n2077), .Y(n1972) );
  NOR2XL U1367 ( .A(work_cntr[14]), .B(n1988), .Y(n1970) );
  NOR4XL U1368 ( .A(n1964), .B(n1963), .C(n1962), .D(n1961), .Y(n1966) );
  NAND3XL U1369 ( .A(n1960), .B(n1959), .C(n1958), .Y(n1961) );
  NAND4XL U1370 ( .A(n1957), .B(n1956), .C(n1955), .D(n1954), .Y(n1962) );
  AOI211XL U1371 ( .A0(n2324), .A1(n2119), .B0(n1953), .C0(n2322), .Y(n1957)
         );
  NAND3XL U1372 ( .A(n1952), .B(n1951), .C(n1950), .Y(n1963) );
  NAND4XL U1373 ( .A(n1949), .B(n1948), .C(n1947), .D(n1946), .Y(n1964) );
  NAND2XL U1374 ( .A(n1943), .B(n1942), .Y(n1944) );
  NAND2XL U1375 ( .A(n1938), .B(n1936), .Y(n1937) );
  INVXL U1376 ( .A(n1940), .Y(n1932) );
  NOR2XL U1377 ( .A(n1939), .B(n1938), .Y(n1930) );
  NAND2XL U1378 ( .A(n1931), .B(n1940), .Y(n1935) );
  NAND2XL U1379 ( .A(n1926), .B(n1925), .Y(n1929) );
  NAND2XL U1380 ( .A(n1921), .B(n1920), .Y(n1925) );
  INVXL U1381 ( .A(n1913), .Y(n1918) );
  NOR2XL U1382 ( .A(n1922), .B(n1912), .Y(n1919) );
  INVXL U1383 ( .A(n1912), .Y(n1924) );
  NOR2XL U1384 ( .A(n1914), .B(n1913), .Y(n1909) );
  NAND2XL U1385 ( .A(n1910), .B(n1915), .Y(n1920) );
  NAND2XL U1386 ( .A(n1905), .B(n1907), .Y(n1915) );
  NAND2XL U1387 ( .A(n121), .B(n1903), .Y(n1907) );
  NAND2XL U1388 ( .A(n1900), .B(n1899), .Y(n1903) );
  NOR2XL U1389 ( .A(n1953), .B(n148), .Y(n1898) );
  INVXL U1390 ( .A(n1947), .Y(n1893) );
  INVXL U1391 ( .A(n148), .Y(n1902) );
  NAND2XL U1392 ( .A(n1892), .B(n1891), .Y(n1900) );
  NAND2XL U1393 ( .A(n1897), .B(n1947), .Y(n1891) );
  NAND2BXL U1394 ( .AN(n1892), .B(n1894), .Y(n1899) );
  NAND2XL U1395 ( .A(n1888), .B(n1890), .Y(n1894) );
  NAND2XL U1396 ( .A(n118), .B(n1886), .Y(n1890) );
  NAND2XL U1397 ( .A(n1884), .B(n1889), .Y(n1883) );
  NOR2XL U1398 ( .A(n1885), .B(n1884), .Y(n1882) );
  INVXL U1399 ( .A(n1948), .Y(n1885) );
  NAND2BXL U1400 ( .AN(n1874), .B(n1878), .Y(n1876) );
  NAND2XL U1401 ( .A(n1873), .B(n1872), .Y(n1878) );
  NAND2XL U1402 ( .A(n1874), .B(n1871), .Y(n1875) );
  NAND2XL U1403 ( .A(n1881), .B(n1956), .Y(n1871) );
  NAND2XL U1404 ( .A(n1869), .B(n1868), .Y(n1872) );
  NAND2XL U1405 ( .A(n1866), .B(n1870), .Y(n1865) );
  NOR2XL U1406 ( .A(n1867), .B(n1866), .Y(n1864) );
  NAND2BXL U1407 ( .AN(n1856), .B(n1860), .Y(n1858) );
  NAND2XL U1408 ( .A(n1855), .B(n1854), .Y(n1860) );
  NAND2XL U1409 ( .A(n1853), .B(n1856), .Y(n1857) );
  NAND2XL U1410 ( .A(n1850), .B(n1848), .Y(n1849) );
  NAND2XL U1411 ( .A(n1863), .B(n1954), .Y(n1853) );
  NOR2XL U1412 ( .A(n1851), .B(n1850), .Y(n1846) );
  NAND2XL U1413 ( .A(n1847), .B(n1852), .Y(n1854) );
  NAND2XL U1414 ( .A(n120), .B(n1841), .Y(n1845) );
  NAND2XL U1415 ( .A(n1837), .B(n1836), .Y(n1841) );
  NOR2XL U1416 ( .A(n1838), .B(n1834), .Y(n1835) );
  INVXL U1417 ( .A(n1955), .Y(n1838) );
  INVXL U1418 ( .A(n1834), .Y(n1840) );
  NAND2XL U1419 ( .A(n1828), .B(n1827), .Y(n1837) );
  NAND2XL U1420 ( .A(n1833), .B(n1952), .Y(n1828) );
  NAND2BXL U1421 ( .AN(n1827), .B(n1830), .Y(n1836) );
  NAND2XL U1422 ( .A(n1823), .B(n1822), .Y(n1826) );
  NAND2XL U1423 ( .A(n1820), .B(n110), .Y(n1819) );
  INVXL U1424 ( .A(n1811), .Y(n1816) );
  NOR2XL U1425 ( .A(n1821), .B(n1820), .Y(n1817) );
  INVXL U1426 ( .A(n1813), .Y(n1808) );
  INVXL U1427 ( .A(n1960), .Y(n1821) );
  INVXL U1428 ( .A(n1818), .Y(n1822) );
  NOR2XL U1429 ( .A(n1812), .B(n1811), .Y(n1806) );
  INVXL U1430 ( .A(n1951), .Y(n1812) );
  NAND2XL U1431 ( .A(n1807), .B(n1813), .Y(n1810) );
  NAND2XL U1432 ( .A(n1803), .B(n1805), .Y(n1813) );
  NAND2BXL U1433 ( .AN(n1802), .B(n1801), .Y(n1805) );
  NAND2XL U1434 ( .A(n1802), .B(n1795), .Y(n1803) );
  NAND2XL U1435 ( .A(n1800), .B(n1958), .Y(n1795) );
  NOR2XL U1436 ( .A(n219), .B(n953), .Y(n954) );
  NAND2XL U1437 ( .A(n1792), .B(n1790), .Y(n1791) );
  NOR2XL U1438 ( .A(n1794), .B(n1792), .Y(n1788) );
  INVXL U1439 ( .A(n1950), .Y(n1794) );
  NAND2XL U1440 ( .A(n1787), .B(n1793), .Y(n1796) );
  INVXL U1441 ( .A(n1789), .Y(n1793) );
  INVXL U1442 ( .A(n1786), .Y(n1782) );
  NAND3XL U1443 ( .A(work_cntr[19]), .B(n1781), .C(n1959), .Y(n1786) );
  NAND2XL U1444 ( .A(n1606), .B(n1708), .Y(n945) );
  NAND2XL U1445 ( .A(n273), .B(N579), .Y(n338) );
  NAND2XL U1446 ( .A(n273), .B(N581), .Y(n339) );
  NAND2XL U1447 ( .A(n273), .B(n272), .Y(n340) );
  NAND2XL U1448 ( .A(n273), .B(N583), .Y(n341) );
  NAND2XL U1449 ( .A(n273), .B(N584), .Y(n342) );
  NAND2XL U1450 ( .A(n2314), .B(n621), .Y(n343) );
  NAND2XL U1451 ( .A(n273), .B(write_addr[8]), .Y(n344) );
  MXI2XL U1452 ( .A(n612), .B(n244), .S0(n273), .Y(n481) );
  NAND2XL U1453 ( .A(n610), .B(n2314), .Y(n346) );
  NAND2XL U1454 ( .A(n2314), .B(n606), .Y(n350) );
  NAND2XL U1455 ( .A(write_addr[12]), .B(n273), .Y(n351) );
  NAND2XL U1456 ( .A(n273), .B(write_addr[13]), .Y(n353) );
  NAND2BXL U1457 ( .AN(n1766), .B(si_sel), .Y(n332) );
  AOI211XL U1458 ( .A0(n1763), .A1(n2331), .B0(n1762), .C0(n1761), .Y(n1766)
         );
  AOI211XL U1459 ( .A0(n1760), .A1(n1759), .B0(n1758), .C0(n1757), .Y(n1762)
         );
  NOR2XL U1460 ( .A(n1760), .B(n1759), .Y(n1757) );
  NAND2XL U1461 ( .A(N2061), .B(n1738), .Y(n1742) );
  NOR4XL U1462 ( .A(n1753), .B(n1752), .C(n1743), .D(n167), .Y(n1736) );
  INVXL U1463 ( .A(n1745), .Y(n1753) );
  NAND4XL U1464 ( .A(n1744), .B(n1745), .C(n1734), .D(n1733), .Y(n1737) );
  NAND2XL U1465 ( .A(n1743), .B(n2097), .Y(n1733) );
  INVXL U1466 ( .A(n1752), .Y(n1744) );
  OAI211XL U1467 ( .A0(N2062), .A1(n1752), .B0(n1745), .C0(n1729), .Y(n1730)
         );
  NOR2BXL U1468 ( .AN(n1721), .B(n2122), .Y(n1723) );
  AND2XL U1469 ( .A(n1728), .B(n1727), .Y(n1731) );
  INVXL U1470 ( .A(n1719), .Y(n1715) );
  NOR2XL U1471 ( .A(n2122), .B(n1714), .Y(n1718) );
  INVXL U1472 ( .A(n1724), .Y(n1714) );
  INVXL U1473 ( .A(n1701), .Y(n1702) );
  OAI211XL U1474 ( .A0(n1697), .A1(n1696), .B0(n1699), .C0(n1700), .Y(n1698)
         );
  NOR2XL U1475 ( .A(n1707), .B(n1706), .Y(n1704) );
  NOR2XL U1476 ( .A(n1690), .B(n1689), .Y(n1692) );
  INVXL U1477 ( .A(n1700), .Y(n1689) );
  AND2XL U1478 ( .A(n1691), .B(n1699), .Y(n1690) );
  INVXL U1479 ( .A(n1682), .Y(n1684) );
  OAI211XL U1480 ( .A0(n1681), .A1(n1682), .B0(n1675), .C0(n1680), .Y(n1677)
         );
  NAND2XL U1481 ( .A(n1674), .B(n1673), .Y(n1680) );
  INVXL U1482 ( .A(n1670), .Y(n1675) );
  INVXL U1483 ( .A(n1667), .Y(n1668) );
  INVXL U1484 ( .A(n1656), .Y(n1662) );
  INVXL U1485 ( .A(n1648), .Y(n1649) );
  NAND2XL U1486 ( .A(n1651), .B(n1647), .Y(n1652) );
  INVXL U1487 ( .A(n1645), .Y(n1642) );
  INVXL U1488 ( .A(n1635), .Y(n1653) );
  NAND2XL U1489 ( .A(n1630), .B(n1632), .Y(n1635) );
  NAND2XL U1490 ( .A(n1627), .B(n1639), .Y(n1637) );
  INVXL U1491 ( .A(n1631), .Y(n1639) );
  NOR2XL U1492 ( .A(work_cntr[19]), .B(n1619), .Y(n1621) );
  NOR2XL U1493 ( .A(n1618), .B(n1617), .Y(n1623) );
  INVXL U1494 ( .A(n1614), .Y(n1620) );
  NAND2XL U1495 ( .A(n1614), .B(n1615), .Y(n1613) );
  NAND2XL U1496 ( .A(n1610), .B(n183), .Y(n1611) );
  INVXL U1497 ( .A(n1671), .Y(n1610) );
  INVXL U1498 ( .A(n1705), .Y(n1710) );
  AOI222XL U1499 ( .A0(n676), .A1(\C162/DATA3_0 ), .B0(n268), .B1(
        global_cntr[0]), .C0(n269), .C1(N1446), .Y(\im_a[0]_BAR ) );
  AOI222XL U1500 ( .A0(n676), .A1(\C162/DATA3_19 ), .B0(global_cntr[19]), .B1(
        n268), .C0(n269), .C1(N1465), .Y(\im_a[19]_BAR ) );
  INVXL U1501 ( .A(n688), .Y(n666) );
  INVXL U1502 ( .A(n664), .Y(n668) );
  NOR2BXL U1503 ( .AN(curr_photo_addr[19]), .B(n266), .Y(\C1/Z_19 ) );
  AOI211XL U1504 ( .A0(n271), .A1(n592), .B0(n576), .C0(n575), .Y(n577) );
  NOR2XL U1505 ( .A(n647), .B(n582), .Y(n576) );
  AOI211XL U1506 ( .A0(n655), .A1(n652), .B0(n651), .C0(n650), .Y(n653) );
  NOR2XL U1507 ( .A(n654), .B(n647), .Y(n651) );
  OAI211XL U1508 ( .A0(n642), .A1(n571), .B0(n565), .C0(n564), .Y(\C163/Z_1 )
         );
  NAND2XL U1509 ( .A(N580), .B(n568), .Y(n564) );
  AOI22XL U1510 ( .A0(N464), .A1(n567), .B0(N580), .B1(n267), .Y(n565) );
  AOI211XL U1511 ( .A0(\intadd_3/B[0] ), .A1(n1054), .B0(n114), .C0(n1353), 
        .Y(n1064) );
  OAI211XL U1512 ( .A0(n640), .A1(n571), .B0(n570), .C0(n569), .Y(\C163/Z_0 )
         );
  NAND2XL U1513 ( .A(N579), .B(n568), .Y(n569) );
  AOI22XL U1514 ( .A0(n238), .A1(n567), .B0(N579), .B1(n267), .Y(n570) );
  NOR2BXL U1515 ( .AN(curr_photo_addr[0]), .B(n266), .Y(n677) );
  AOI211XL U1516 ( .A0(n645), .A1(n652), .B0(n644), .C0(n643), .Y(n646) );
  NOR2XL U1517 ( .A(n642), .B(n641), .Y(n644) );
  INVXL U1518 ( .A(n640), .Y(n652) );
  NOR2XL U1519 ( .A(n1355), .B(N579), .Y(n337) );
  AOI211XL U1520 ( .A0(\intadd_3/A[0] ), .A1(n1201), .B0(n1353), .C0(n1200), 
        .Y(n1202) );
  NOR2XL U1521 ( .A(\intadd_3/A[0] ), .B(n1201), .Y(n1200) );
  OAI211XL U1522 ( .A0(n563), .A1(n162), .B0(n562), .C0(n561), .Y(\C163/Z_2 )
         );
  NAND2XL U1523 ( .A(n1372), .B(n638), .Y(n561) );
  AOI22XL U1524 ( .A0(N465), .A1(n567), .B0(N581), .B1(n267), .Y(n562) );
  AOI211XL U1525 ( .A0(n655), .A1(n638), .B0(n637), .C0(n636), .Y(n639) );
  NOR2XL U1526 ( .A(n642), .B(n647), .Y(n637) );
  OAI211XL U1527 ( .A0(n632), .A1(n571), .B0(n560), .C0(n559), .Y(\C163/Z_3 )
         );
  NAND2XL U1528 ( .A(n272), .B(n568), .Y(n559) );
  AOI22XL U1529 ( .A0(N466), .A1(n567), .B0(n272), .B1(n267), .Y(n560) );
  AOI211XL U1530 ( .A0(n645), .A1(n638), .B0(n634), .C0(n633), .Y(n635) );
  NOR2XL U1531 ( .A(n632), .B(n641), .Y(n634) );
  OAI211XL U1532 ( .A0(n563), .A1(n2310), .B0(n558), .C0(n557), .Y(\C163/Z_4 )
         );
  NAND2XL U1533 ( .A(n1372), .B(n629), .Y(n557) );
  AOI22XL U1534 ( .A0(N467), .A1(n567), .B0(N583), .B1(n267), .Y(n558) );
  NOR2BXL U1535 ( .AN(curr_photo_addr[5]), .B(n266), .Y(\C1/Z_5 ) );
  AOI211XL U1536 ( .A0(n655), .A1(n629), .B0(n628), .C0(n627), .Y(n631) );
  NOR2XL U1537 ( .A(n632), .B(n647), .Y(n628) );
  OAI211XL U1538 ( .A0(n1348), .A1(n272), .B0(n718), .C0(n1347), .Y(n1349) );
  OAI211XL U1539 ( .A0(n623), .A1(n571), .B0(n556), .C0(n555), .Y(\C163/Z_5 )
         );
  NAND2XL U1540 ( .A(N584), .B(n568), .Y(n555) );
  AOI22XL U1541 ( .A0(N468), .A1(n567), .B0(N584), .B1(n267), .Y(n556) );
  NOR2BXL U1542 ( .AN(curr_photo_addr[6]), .B(n266), .Y(\C1/Z_6 ) );
  AOI211XL U1543 ( .A0(n645), .A1(n629), .B0(n625), .C0(n624), .Y(n626) );
  NOR2XL U1544 ( .A(n623), .B(n641), .Y(n625) );
  OAI211XL U1545 ( .A0(n563), .A1(n241), .B0(n554), .C0(n553), .Y(\C163/Z_6 )
         );
  NAND2XL U1546 ( .A(n1372), .B(n621), .Y(n553) );
  AOI22XL U1547 ( .A0(N469), .A1(n567), .B0(N585), .B1(n267), .Y(n554) );
  AOI211XL U1548 ( .A0(n655), .A1(n621), .B0(n620), .C0(n619), .Y(n622) );
  NOR2XL U1549 ( .A(n623), .B(n647), .Y(n620) );
  OAI211XL U1550 ( .A0(n612), .A1(n571), .B0(n552), .C0(n551), .Y(\C163/Z_7 )
         );
  NAND2XL U1551 ( .A(write_addr[9]), .B(n568), .Y(n551) );
  AOI22XL U1552 ( .A0(N470), .A1(n567), .B0(n244), .B1(n267), .Y(n552) );
  NOR2BXL U1553 ( .AN(curr_photo_addr[8]), .B(n266), .Y(\C1/Z_8 ) );
  AOI211XL U1554 ( .A0(n645), .A1(n621), .B0(n617), .C0(n616), .Y(n618) );
  NOR2XL U1555 ( .A(n615), .B(n641), .Y(n617) );
  OAI211XL U1556 ( .A0(n563), .A1(n243), .B0(n550), .C0(n549), .Y(\C163/Z_8 )
         );
  NAND2XL U1557 ( .A(n1372), .B(n610), .Y(n549) );
  AOI22XL U1558 ( .A0(N471), .A1(n567), .B0(N587), .B1(n267), .Y(n550) );
  NOR2BXL U1559 ( .AN(curr_photo_addr[9]), .B(n266), .Y(\C1/Z_9 ) );
  INVXL U1560 ( .A(n660), .Y(n614) );
  OAI211XL U1561 ( .A0(n563), .A1(n245), .B0(n548), .C0(n547), .Y(\C163/Z_9 )
         );
  NAND2XL U1562 ( .A(n1372), .B(n606), .Y(n547) );
  AOI22XL U1563 ( .A0(N472), .A1(n567), .B0(N588), .B1(n267), .Y(n548) );
  NOR2BXL U1564 ( .AN(curr_photo_addr[10]), .B(n266), .Y(\C1/Z_10 ) );
  AOI211XL U1565 ( .A0(n655), .A1(n610), .B0(n609), .C0(n608), .Y(n611) );
  NOR2XL U1566 ( .A(n615), .B(n647), .Y(n609) );
  AOI211XL U1567 ( .A0(n1330), .A1(n1297), .B0(n2284), .C0(n1245), .Y(n1246)
         );
  OAI211XL U1568 ( .A0(n563), .A1(n164), .B0(n546), .C0(n545), .Y(\C163/Z_10 )
         );
  NAND2XL U1569 ( .A(n1372), .B(n595), .Y(n545) );
  AOI22XL U1570 ( .A0(N473), .A1(n567), .B0(N589), .B1(n267), .Y(n546) );
  AOI211XL U1571 ( .A0(n655), .A1(n606), .B0(n605), .C0(n604), .Y(n607) );
  NOR2XL U1572 ( .A(n612), .B(n647), .Y(n605) );
  NOR2BXL U1573 ( .AN(curr_photo_addr[12]), .B(n266), .Y(\C1/Z_12 ) );
  AOI211XL U1574 ( .A0(n645), .A1(n610), .B0(n602), .C0(n601), .Y(n603) );
  NOR2XL U1575 ( .A(n600), .B(n641), .Y(n602) );
  INVXL U1576 ( .A(n595), .Y(n600) );
  AOI211XL U1577 ( .A0(n1242), .A1(n1243), .B0(n1289), .C0(n1327), .Y(n1244)
         );
  INVXL U1578 ( .A(n1296), .Y(n1242) );
  OAI211XL U1579 ( .A0(n594), .A1(n571), .B0(n544), .C0(n543), .Y(\C163/Z_12 )
         );
  NAND2XL U1580 ( .A(write_addr[14]), .B(n568), .Y(n543) );
  AOI22XL U1581 ( .A0(N475), .A1(n567), .B0(N591), .B1(n267), .Y(n544) );
  AOI211XL U1582 ( .A0(n645), .A1(n606), .B0(n598), .C0(n597), .Y(n599) );
  NOR2XL U1583 ( .A(n596), .B(n641), .Y(n598) );
  AOI211XL U1584 ( .A0(write_addr[11]), .A1(n348), .B0(n1293), .C0(n347), .Y(
        n349) );
  NOR2XL U1585 ( .A(n1355), .B(n1292), .Y(n347) );
  AOI211XL U1586 ( .A0(n1292), .A1(n1291), .B0(n1290), .C0(n1327), .Y(n1293)
         );
  INVXL U1587 ( .A(n1303), .Y(n1290) );
  INVXL U1588 ( .A(n265), .Y(n348) );
  XOR2XL U1589 ( .A(\intadd_4/A[2] ), .B(\intadd_4/n3 ), .Y(\intadd_4/SUM[2] )
         );
  OAI211XL U1590 ( .A0(n108), .A1(n571), .B0(n542), .C0(n541), .Y(\C163/Z_13 )
         );
  NAND2XL U1591 ( .A(write_addr[15]), .B(n568), .Y(n541) );
  AOI22XL U1592 ( .A0(N476), .A1(n567), .B0(N592), .B1(n267), .Y(n542) );
  AOI211XL U1593 ( .A0(n1304), .A1(n1303), .B0(n1311), .C0(n1327), .Y(n1305)
         );
  XOR2XL U1594 ( .A(\intadd_4/B[3] ), .B(n191), .Y(\intadd_4/SUM[3] ) );
  AOI211XL U1595 ( .A0(write_addr[13]), .A1(n592), .B0(n591), .C0(n590), .Y(
        n593) );
  NOR2XL U1596 ( .A(n596), .B(n647), .Y(n591) );
  NOR2XL U1597 ( .A(n265), .B(n166), .Y(n352) );
  AOI211XL U1598 ( .A0(n1323), .A1(n1322), .B0(n1308), .C0(n1307), .Y(n1309)
         );
  NOR2XL U1599 ( .A(n1323), .B(n1322), .Y(n1307) );
  AND2XL U1600 ( .A(\intadd_4/B[3] ), .B(n191), .Y(n192) );
  AND2XL U1601 ( .A(\intadd_4/A[2] ), .B(\intadd_4/n3 ), .Y(n191) );
  INVXL U1602 ( .A(\intadd_3/n1 ), .Y(\intadd_4/B[1] ) );
  INVXL U1603 ( .A(n1219), .Y(\intadd_3/B[1] ) );
  INVXL U1604 ( .A(n1216), .Y(\intadd_3/A[1] ) );
  AOI21XL U1605 ( .A0(n1229), .A1(n1215), .B0(n1221), .Y(n1342) );
  NAND2XL U1606 ( .A(n1209), .B(n1208), .Y(n1210) );
  NOR2XL U1607 ( .A(n1209), .B(n1208), .Y(n1211) );
  INVXL U1608 ( .A(n1206), .Y(n1197) );
  NAND2XL U1609 ( .A(n1773), .B(\next_cr_y[0] ), .Y(n1198) );
  INVXL U1610 ( .A(n1196), .Y(n1773) );
  INVXL U1611 ( .A(\intadd_3/SUM[0] ), .Y(n1344) );
  NAND2XL U1612 ( .A(n1207), .B(n1224), .Y(\intadd_3/CI ) );
  NAND2BXL U1613 ( .AN(n1049), .B(n1048), .Y(n1050) );
  AOI211XL U1614 ( .A0(\intadd_3/A[0] ), .A1(n1771), .B0(n1042), .C0(n1041), 
        .Y(n1043) );
  NOR2XL U1615 ( .A(n1027), .B(n1224), .Y(n1037) );
  NAND2BXL U1616 ( .AN(n1031), .B(n1049), .Y(n1047) );
  INVXL U1617 ( .A(n1225), .Y(\intadd_3/B[2] ) );
  INVXL U1618 ( .A(n1222), .Y(\intadd_3/A[2] ) );
  AND2XL U1619 ( .A(n1203), .B(\next_cr_y[0] ), .Y(n1213) );
  INVXL U1620 ( .A(n1232), .Y(\intadd_3/B[3] ) );
  INVXL U1621 ( .A(n1228), .Y(\intadd_3/A[3] ) );
  INVXL U1622 ( .A(n1032), .Y(n1035) );
  AND3XL U1623 ( .A(n1030), .B(n1028), .C(n1224), .Y(n1021) );
  NAND2XL U1624 ( .A(n1028), .B(n1224), .Y(n1029) );
  INVXL U1625 ( .A(n1236), .Y(\intadd_3/B[4] ) );
  INVXL U1626 ( .A(n1235), .Y(\intadd_3/A[4] ) );
  INVXL U1627 ( .A(n1016), .Y(n1019) );
  NAND2XL U1628 ( .A(n1020), .B(n1034), .Y(n1033) );
  AND3XL U1629 ( .A(n1012), .B(n1011), .C(n1231), .Y(n1014) );
  NAND3XL U1630 ( .A(n1022), .B(n1030), .C(n1028), .Y(n1020) );
  NAND2XL U1631 ( .A(n1231), .B(n1023), .Y(n1024) );
  INVXL U1632 ( .A(n1239), .Y(\intadd_3/B[5] ) );
  INVXL U1633 ( .A(n1003), .Y(n1006) );
  NAND2XL U1634 ( .A(n1018), .B(n1013), .Y(n1017) );
  NAND3XL U1635 ( .A(n1012), .B(n1015), .C(n1011), .Y(n1013) );
  NAND2XL U1636 ( .A(n1002), .B(n1237), .Y(n1008) );
  NOR2XL U1637 ( .A(n994), .B(next_cr_x[5]), .Y(n996) );
  AND3XL U1638 ( .A(n1001), .B(n999), .C(n1237), .Y(n992) );
  INVXL U1639 ( .A(n968), .Y(n971) );
  NAND2XL U1640 ( .A(n1005), .B(n991), .Y(n1004) );
  NAND3XL U1641 ( .A(n1001), .B(n993), .C(n999), .Y(n991) );
  NOR2BXL U1642 ( .AN(n965), .B(n1223), .Y(n959) );
  NAND2XL U1643 ( .A(n994), .B(next_cr_x[5]), .Y(n995) );
  NOR2XL U1644 ( .A(n961), .B(next_cr_x[6]), .Y(n962) );
  XNOR2XL U1645 ( .A(n262), .B(next_cr_x[6]), .Y(n207) );
  XOR2XL U1646 ( .A(\next_cr_y[0] ), .B(next_cr_x[5]), .Y(n262) );
  INVXL U1647 ( .A(\intadd_4/SUM[0] ), .Y(\intadd_3/B[6] ) );
  MX2XL U1648 ( .A(n263), .B(n264), .S0(next_cr_x[5]), .Y(n206) );
  NAND2XL U1649 ( .A(n970), .B(n958), .Y(n969) );
  NAND2XL U1650 ( .A(n960), .B(n965), .Y(n958) );
  NOR2BXL U1651 ( .AN(n764), .B(n1230), .Y(n765) );
  AND3XL U1652 ( .A(n764), .B(n175), .C(next_cr_x[6]), .Y(n762) );
  NAND2BXL U1653 ( .AN(\next_cr_y[0] ), .B(next_cr_x[6]), .Y(n264) );
  NAND2XL U1654 ( .A(next_cr_x[6]), .B(\next_cr_y[0] ), .Y(n263) );
  NAND2XL U1655 ( .A(n1203), .B(n1214), .Y(n1212) );
  INVXL U1656 ( .A(n901), .Y(n905) );
  NOR2XL U1657 ( .A(n1288), .B(n898), .Y(n899) );
  INVXL U1658 ( .A(n897), .Y(n903) );
  AOI211XL U1659 ( .A0(n224), .A1(n185), .B0(n270), .C0(n882), .Y(n772) );
  NAND3XL U1660 ( .A(n763), .B(n764), .C(n175), .Y(n761) );
  NAND2XL U1661 ( .A(n769), .B(n768), .Y(n764) );
  INVXL U1662 ( .A(n786), .Y(n763) );
  INVXL U1663 ( .A(n1288), .Y(\intadd_4/A[1] ) );
  NAND3XL U1664 ( .A(n892), .B(n1301), .C(n891), .Y(n890) );
  NOR2XL U1665 ( .A(n895), .B(n896), .Y(n893) );
  NOR2XL U1666 ( .A(n1287), .B(n1040), .Y(n888) );
  NAND2XL U1667 ( .A(n887), .B(n886), .Y(n889) );
  NAND2XL U1668 ( .A(n1299), .B(n1287), .Y(n1286) );
  NAND3XL U1669 ( .A(n1302), .B(n1299), .C(n1301), .Y(n1300) );
  NAND3XL U1670 ( .A(n1285), .B(n1281), .C(n1284), .Y(n1282) );
  NAND2XL U1671 ( .A(n874), .B(n875), .Y(n873) );
  INVXL U1672 ( .A(n872), .Y(n875) );
  NOR2BXL U1673 ( .AN(n892), .B(n891), .Y(n876) );
  INVXL U1674 ( .A(n866), .Y(n870) );
  INVXL U1675 ( .A(n868), .Y(n871) );
  NAND3XL U1676 ( .A(n865), .B(n867), .C(n1771), .Y(n863) );
  NOR2BXL U1677 ( .AN(n1771), .B(n1285), .Y(n864) );
  INVXL U1678 ( .A(n877), .Y(n880) );
  NAND2XL U1679 ( .A(n1774), .B(n887), .Y(n877) );
  INVXL U1680 ( .A(n1298), .Y(n1302) );
  NAND3XL U1681 ( .A(n1283), .B(n1278), .C(n1280), .Y(n1279) );
  NAND2XL U1682 ( .A(n1284), .B(n1281), .Y(n1278) );
  NAND2XL U1683 ( .A(n1277), .B(n1276), .Y(n1281) );
  NAND3XL U1684 ( .A(n113), .B(n1277), .C(n860), .Y(n859) );
  NOR2XL U1685 ( .A(n874), .B(n872), .Y(n862) );
  NOR2XL U1686 ( .A(n1274), .B(n1027), .Y(n852) );
  NAND2XL U1687 ( .A(n851), .B(n854), .Y(n853) );
  NAND2XL U1688 ( .A(n1277), .B(n1275), .Y(n1273) );
  NOR2BXL U1689 ( .AN(n113), .B(n860), .Y(n850) );
  INVXL U1690 ( .A(n843), .Y(n857) );
  NAND2XL U1691 ( .A(n841), .B(n839), .Y(n840) );
  NAND2XL U1692 ( .A(n1776), .B(n1269), .Y(n839) );
  INVXL U1693 ( .A(n855), .Y(n858) );
  NAND2XL U1694 ( .A(n1775), .B(n851), .Y(n855) );
  INVXL U1695 ( .A(n775), .Y(n778) );
  NAND2XL U1696 ( .A(n1270), .B(n1269), .Y(n1271) );
  INVXL U1697 ( .A(n846), .Y(n842) );
  NAND2XL U1698 ( .A(n837), .B(n838), .Y(n836) );
  INVXL U1699 ( .A(n835), .Y(n838) );
  OAI31XL U1700 ( .A0(n834), .A1(n833), .A2(n832), .B0(n831), .Y(n849) );
  INVXL U1701 ( .A(n830), .Y(n832) );
  INVXL U1702 ( .A(n829), .Y(n834) );
  INVXL U1703 ( .A(n1264), .Y(n1266) );
  NOR2XL U1704 ( .A(n1261), .B(n1263), .Y(n1260) );
  NAND2XL U1705 ( .A(n1256), .B(n1255), .Y(n1258) );
  NOR2XL U1706 ( .A(n1251), .B(n184), .Y(n1253) );
  NAND2XL U1707 ( .A(n184), .B(n1251), .Y(n1250) );
  NAND2XL U1708 ( .A(n825), .B(n824), .Y(n826) );
  NOR2XL U1709 ( .A(n835), .B(n837), .Y(n827) );
  NAND2XL U1710 ( .A(n828), .B(n1778), .Y(n829) );
  INVXL U1711 ( .A(n779), .Y(n782) );
  NAND2XL U1712 ( .A(n822), .B(n820), .Y(n821) );
  NAND2XL U1713 ( .A(n115), .B(n1256), .Y(n820) );
  INVXL U1714 ( .A(n816), .Y(n823) );
  NAND2XL U1715 ( .A(n813), .B(n814), .Y(n812) );
  INVXL U1716 ( .A(n811), .Y(n814) );
  NOR2BXL U1717 ( .AN(n824), .B(n825), .Y(n815) );
  NAND2BXL U1718 ( .AN(n813), .B(n1252), .Y(n809) );
  NAND3XL U1719 ( .A(n806), .B(n810), .C(n1779), .Y(n804) );
  NOR2XL U1720 ( .A(n1251), .B(n961), .Y(n805) );
  NAND3XL U1721 ( .A(n802), .B(n1249), .C(n801), .Y(n800) );
  NOR2XL U1722 ( .A(n813), .B(n811), .Y(n803) );
  INVXL U1723 ( .A(n795), .Y(n796) );
  NAND2XL U1724 ( .A(n1779), .B(n806), .Y(n808) );
  NAND2XL U1725 ( .A(n790), .B(n771), .Y(n789) );
  NOR2BXL U1726 ( .AN(n802), .B(n801), .Y(n791) );
  INVXL U1727 ( .A(n787), .Y(n786) );
  INVXL U1728 ( .A(n785), .Y(n788) );
  INVXL U1729 ( .A(n175), .Y(n261) );
  NAND2XL U1730 ( .A(n1780), .B(n175), .Y(n785) );
  INVXL U1731 ( .A(n964), .Y(n792) );
  AOI211XL U1732 ( .A0(n107), .A1(n759), .B0(n757), .C0(n270), .Y(n758) );
  OAI211XL U1733 ( .A0(write_cntr[9]), .A1(n766), .B0(n759), .C0(n783), .Y(
        n760) );
  NOR2XL U1734 ( .A(n2288), .B(n2289), .Y(n884) );
  INVXL U1735 ( .A(n750), .Y(n1761) );
  INVXL U1736 ( .A(n748), .Y(n749) );
  NOR3XL U1737 ( .A(n1777), .B(n209), .C(n173), .Y(n747) );
  NAND2XL U1738 ( .A(write_cntr[6]), .B(n780), .Y(n779) );
  NAND2XL U1739 ( .A(n776), .B(write_cntr[4]), .Y(n775) );
  OAI211XL U1740 ( .A0(n582), .A1(n571), .B0(n540), .C0(n539), .Y(\C163/Z_15 )
         );
  NAND2XL U1741 ( .A(n271), .B(n568), .Y(n539) );
  AOI22XL U1742 ( .A0(N478), .A1(n567), .B0(N594), .B1(n267), .Y(n540) );
  NOR2BXL U1743 ( .AN(curr_photo_addr[16]), .B(n266), .Y(\C1/Z_16 ) );
  AOI211XL U1744 ( .A0(write_addr[14]), .A1(n592), .B0(n588), .C0(n587), .Y(
        n589) );
  NOR2XL U1745 ( .A(n594), .B(n647), .Y(n588) );
  AOI211XL U1746 ( .A0(n1312), .A1(n1317), .B0(n1318), .C0(n1327), .Y(n1313)
         );
  INVXL U1747 ( .A(n1312), .Y(n334) );
  OAI211XL U1748 ( .A0(n2313), .A1(n571), .B0(n538), .C0(n533), .Y(\C163/Z_16 ) );
  NAND2XL U1749 ( .A(write_addr[18]), .B(n521), .Y(n533) );
  AOI22XL U1750 ( .A0(N479), .A1(n567), .B0(N595), .B1(n267), .Y(n538) );
  NOR2BXL U1751 ( .AN(curr_photo_addr[17]), .B(n266), .Y(\C1/Z_17 ) );
  AOI211XL U1752 ( .A0(write_addr[15]), .A1(n592), .B0(n584), .C0(n583), .Y(
        n585) );
  NOR2XL U1753 ( .A(n108), .B(n647), .Y(n584) );
  NAND2XL U1754 ( .A(write_addr[14]), .B(n1314), .Y(n1316) );
  INVXL U1755 ( .A(n1310), .Y(n1314) );
  OAI211XL U1756 ( .A0(n574), .A1(n571), .B0(n520), .C0(n517), .Y(\C163/Z_17 )
         );
  NAND2XL U1757 ( .A(write_addr[19]), .B(n521), .Y(n517) );
  AOI211XL U1758 ( .A0(n1361), .A1(n510), .B0(n170), .C0(n1968), .Y(n511) );
  INVXL U1759 ( .A(n685), .Y(n510) );
  INVXL U1760 ( .A(n1368), .Y(n516) );
  AOI22XL U1761 ( .A0(n112), .A1(n567), .B0(N596), .B1(n267), .Y(n520) );
  OAI211XL U1762 ( .A0(n1364), .A1(n170), .B0(n691), .C0(n1363), .Y(n1367) );
  NAND2XL U1763 ( .A(n1605), .B(n1364), .Y(n1363) );
  NAND2XL U1764 ( .A(n1968), .B(n165), .Y(n1369) );
  INVXL U1765 ( .A(n1333), .Y(n1335) );
  NOR2BXL U1766 ( .AN(curr_photo_addr[18]), .B(n266), .Y(\C1/Z_18 ) );
  AOI211XL U1767 ( .A0(write_addr[16]), .A1(n592), .B0(n580), .C0(n579), .Y(
        n581) );
  INVXL U1768 ( .A(n151), .Y(n1332) );
  INVXL U1769 ( .A(n648), .Y(n656) );
  NOR2XL U1770 ( .A(n586), .B(n647), .Y(n580) );
  NOR2XL U1771 ( .A(n265), .B(n248), .Y(n354) );
  NAND2BXL U1772 ( .AN(n277), .B(n2281), .Y(n1352) );
  NOR2XL U1773 ( .A(n1308), .B(n2), .Y(n355) );
  INVXL U1774 ( .A(n1291), .Y(n1289) );
  NAND2XL U1775 ( .A(write_addr[10]), .B(n1296), .Y(n1291) );
  AOI211XL U1776 ( .A0(n272), .A1(n1346), .B0(n1350), .C0(n1351), .Y(n989) );
  NOR4XL U1777 ( .A(n1334), .B(n1328), .C(n1326), .D(n985), .Y(n990) );
  AOI211XL U1778 ( .A0(n1292), .A1(n1304), .B0(n1358), .C0(n1323), .Y(n985) );
  AND2XL U1779 ( .A(n1315), .B(write_addr[16]), .Y(n981) );
  INVXL U1780 ( .A(n1241), .Y(n982) );
  NAND2XL U1781 ( .A(n1294), .B(write_addr[10]), .Y(n1241) );
  NAND2BXL U1782 ( .AN(n746), .B(n1060), .Y(next_state[1]) );
  INVX6 U1783 ( .A(n2340), .Y(n277) );
  NOR2X2 U1784 ( .A(n746), .B(n2280), .Y(n14) );
  OAI21X1 U1785 ( .A0(n172), .A1(n742), .B0(n743), .Y(n2280) );
  AOI211XL U1786 ( .A0(n2279), .A1(n1516), .B0(n171), .C0(en_so), .Y(n741) );
  NAND3X1 U1787 ( .A(write_cntr[14]), .B(write_cntr[11]), .C(n720), .Y(n721)
         );
  INVXL U1788 ( .A(n739), .Y(n2316) );
  NAND2XL U1789 ( .A(n708), .B(n2279), .Y(n739) );
  NAND4XL U1790 ( .A(n735), .B(n734), .C(n733), .D(n732), .Y(n736) );
  NOR4XL U1791 ( .A(n694), .B(n700), .C(n699), .D(n701), .Y(n732) );
  INVXL U1792 ( .A(n288), .Y(n289) );
  NOR4XL U1793 ( .A(n702), .B(n705), .C(n706), .D(n707), .Y(n733) );
  AOI21X1 U1794 ( .A0(n190), .A1(n280), .B0(n281), .Y(n706) );
  INVXL U1795 ( .A(n738), .Y(n298) );
  NAND2BXL U1796 ( .AN(n731), .B(n728), .Y(n727) );
  NAND2X1 U1797 ( .A(global_cntr[18]), .B(n297), .Y(n728) );
  AOI21X1 U1798 ( .A0(n199), .A1(n294), .B0(n295), .Y(n695) );
  INVXL U1799 ( .A(n294), .Y(n292) );
  AOI21X1 U1800 ( .A0(n198), .A1(n290), .B0(n291), .Y(n698) );
  NOR2X1 U1801 ( .A(n290), .B(n198), .Y(n291) );
  OAI21X1 U1802 ( .A0(global_cntr[9]), .A1(n285), .B0(n286), .Y(n730) );
  AOI21X1 U1803 ( .A0(n194), .A1(n283), .B0(n284), .Y(n703) );
  NOR2XL U1804 ( .A(n726), .B(n729), .Y(n282) );
  NAND2XL U1805 ( .A(n723), .B(n722), .Y(n1514) );
  INVXL U1806 ( .A(n286), .Y(n287) );
  NAND3X1 U1807 ( .A(n284), .B(global_cntr[9]), .C(global_cntr[8]), .Y(n286)
         );
  NOR2X2 U1808 ( .A(n283), .B(n194), .Y(n284) );
  NAND2X1 U1809 ( .A(n708), .B(global_cntr[3]), .Y(n280) );
  INVXL U1810 ( .A(n2330), .Y(n657) );
  NOR2BXL U1811 ( .AN(n684), .B(n1763), .Y(n361) );
  NAND2XL U1812 ( .A(n1192), .B(n1939), .Y(n1193) );
  INVXL U1813 ( .A(n1191), .Y(n1192) );
  INVXL U1814 ( .A(n681), .Y(n573) );
  NAND2XL U1815 ( .A(en_so), .B(n367), .Y(n368) );
  NAND2XL U1816 ( .A(n685), .B(n1511), .Y(n1371) );
  NOR3XL U1817 ( .A(n509), .B(write_addr[8]), .C(n685), .Y(n507) );
  NAND2XL U1818 ( .A(n691), .B(read_cntr[0]), .Y(n509) );
  NAND2XL U1819 ( .A(read_cntr[1]), .B(n1511), .Y(n505) );
  NOR4XL U1820 ( .A(n271), .B(write_addr[16]), .C(write_addr[18]), .D(n166), 
        .Y(n1359) );
  NOR4XL U1821 ( .A(write_addr[19]), .B(n1358), .C(n165), .D(n1357), .Y(n1360)
         );
  NAND2XL U1822 ( .A(n988), .B(N585), .Y(n1356) );
  INVX4 U1823 ( .A(n2334), .Y(si_sel) );
  NAND2XL U1824 ( .A(n667), .B(n688), .Y(n330) );
  NOR2XL U1825 ( .A(n369), .B(n663), .Y(n328) );
  NAND2BXL U1826 ( .AN(n1510), .B(n327), .Y(n667) );
  NOR2XL U1827 ( .A(n2321), .B(n2327), .Y(n1510) );
  INVXL U1828 ( .A(n1188), .Y(n1186) );
  INVXL U1829 ( .A(n1173), .Y(n1175) );
  INVXL U1830 ( .A(n1170), .Y(n1172) );
  INVXL U1831 ( .A(n1181), .Y(n1180) );
  AOI21XL U1832 ( .A0(n1177), .A1(n1173), .B0(n1174), .Y(n1169) );
  NAND2XL U1833 ( .A(n1166), .B(n1171), .Y(n1165) );
  INVXL U1834 ( .A(n1162), .Y(n1160) );
  NOR2XL U1835 ( .A(work_cntr[4]), .B(n1164), .Y(n1157) );
  INVXL U1836 ( .A(n1158), .Y(n1151) );
  NAND2XL U1837 ( .A(n2057), .B(n1163), .Y(n1156) );
  NAND2XL U1838 ( .A(n1687), .B(n1163), .Y(n1136) );
  INVXL U1839 ( .A(n1144), .Y(n1145) );
  INVXL U1840 ( .A(n1148), .Y(n1134) );
  NAND2XL U1841 ( .A(n1135), .B(n226), .Y(n1128) );
  NAND3XL U1842 ( .A(n1126), .B(n1137), .C(n1138), .Y(n1131) );
  NAND2BXL U1843 ( .AN(n1125), .B(n1124), .Y(n1138) );
  NAND2XL U1844 ( .A(n1123), .B(n1125), .Y(n1137) );
  NAND2BXL U1845 ( .AN(n1124), .B(n1118), .Y(n1126) );
  NAND2XL U1846 ( .A(n1120), .B(n1119), .Y(n1124) );
  NOR3XL U1847 ( .A(n1116), .B(n1115), .C(n1114), .Y(n1117) );
  INVXL U1848 ( .A(n1123), .Y(n1118) );
  INVXL U1849 ( .A(n1108), .Y(n1116) );
  NAND2XL U1850 ( .A(n1127), .B(n183), .Y(n1103) );
  INVXL U1851 ( .A(n1112), .Y(n1113) );
  INVXL U1852 ( .A(n1114), .Y(n1101) );
  NAND3XL U1853 ( .A(n1105), .B(n1095), .C(n1104), .Y(n1099) );
  NAND2XL U1854 ( .A(n1094), .B(n1093), .Y(n1104) );
  AND3XL U1855 ( .A(n1127), .B(n183), .C(n222), .Y(n1102) );
  NAND3XL U1856 ( .A(n1092), .B(n1088), .C(n1089), .Y(n1095) );
  NAND2XL U1857 ( .A(n1087), .B(n1086), .Y(n1089) );
  INVXL U1858 ( .A(n1088), .Y(n1094) );
  NAND2BXL U1859 ( .AN(n1079), .B(n1081), .Y(n1082) );
  NAND2XL U1860 ( .A(n1074), .B(n1073), .Y(n1071) );
  NAND2XL U1861 ( .A(work_cntr[19]), .B(n1068), .Y(n1069) );
  NOR2BXL U1862 ( .AN(n1066), .B(work_cntr[17]), .Y(n1067) );
  NAND2XL U1863 ( .A(n1078), .B(n219), .Y(n1077) );
  INVXL U1864 ( .A(n1911), .Y(n1914) );
  NAND2XL U1865 ( .A(n1975), .B(n1163), .Y(n1068) );
  NOR2XL U1866 ( .A(n167), .B(n2331), .Y(n957) );
  NAND2X2 U1867 ( .A(N2061), .B(N85), .Y(n2331) );
  NOR2X2 U1868 ( .A(state[0]), .B(n2328), .Y(n691) );
  NOR2X1 U1869 ( .A(N2062), .B(N2063), .Y(n1374) );
  INVXL U1870 ( .A(n1739), .Y(n326) );
  NAND2BXL U1871 ( .AN(n1507), .B(n324), .Y(n669) );
  NAND2XL U1872 ( .A(n1508), .B(n1509), .Y(n324) );
  NAND2XL U1873 ( .A(n1498), .B(n1497), .Y(n1502) );
  INVXL U1874 ( .A(n1501), .Y(n1503) );
  INVXL U1875 ( .A(n1496), .Y(n1500) );
  NAND2XL U1876 ( .A(n1495), .B(n1496), .Y(n1501) );
  NAND2XL U1877 ( .A(n1492), .B(n1494), .Y(n1496) );
  NAND2XL U1878 ( .A(n119), .B(n1490), .Y(n1494) );
  NAND2XL U1879 ( .A(n1487), .B(n1486), .Y(n1490) );
  NOR2XL U1880 ( .A(N2062), .B(n1484), .Y(n1485) );
  INVXL U1881 ( .A(n1484), .Y(n1489) );
  NAND2XL U1882 ( .A(n1479), .B(n1478), .Y(n1487) );
  NAND2XL U1883 ( .A(n1483), .B(n179), .Y(n1478) );
  NAND2BXL U1884 ( .AN(n1479), .B(n1480), .Y(n1486) );
  NAND2XL U1885 ( .A(n1475), .B(n1477), .Y(n1480) );
  NAND2XL U1886 ( .A(n1474), .B(n1473), .Y(n1477) );
  NAND2XL U1887 ( .A(n1472), .B(n1476), .Y(n1471) );
  NOR2XL U1888 ( .A(work_cntr[4]), .B(n1472), .Y(n1470) );
  NAND2BXL U1889 ( .AN(n1463), .B(n1466), .Y(n1465) );
  NAND2XL U1890 ( .A(n1463), .B(n1460), .Y(n1464) );
  NAND2XL U1891 ( .A(n1469), .B(n168), .Y(n1460) );
  NAND2XL U1892 ( .A(n1458), .B(n1457), .Y(n1461) );
  NAND2XL U1893 ( .A(n1456), .B(n1459), .Y(n1455) );
  NOR2XL U1894 ( .A(work_cntr[6]), .B(n1456), .Y(n1453) );
  INVXL U1895 ( .A(n1449), .Y(n1446) );
  INVXL U1896 ( .A(n1454), .Y(n1457) );
  NAND2XL U1897 ( .A(n1452), .B(n176), .Y(n1445) );
  NAND2XL U1898 ( .A(n1444), .B(n1449), .Y(n1448) );
  NAND2XL U1899 ( .A(n1441), .B(n1443), .Y(n1449) );
  NAND2BXL U1900 ( .AN(n1440), .B(n1439), .Y(n1443) );
  NAND2XL U1901 ( .A(n1437), .B(n1436), .Y(n1439) );
  NAND2BXL U1902 ( .AN(n1432), .B(n1433), .Y(n1436) );
  NAND2BXL U1903 ( .AN(n1429), .B(n1431), .Y(n1433) );
  NAND2XL U1904 ( .A(n1428), .B(n1427), .Y(n1431) );
  NAND2XL U1905 ( .A(n1426), .B(n1430), .Y(n1425) );
  INVXL U1906 ( .A(n1427), .Y(n1424) );
  INVXL U1907 ( .A(n1418), .Y(n1422) );
  NOR2XL U1908 ( .A(work_cntr[10]), .B(n1426), .Y(n1423) );
  NAND2XL U1909 ( .A(n122), .B(n1419), .Y(n1417) );
  NAND2XL U1910 ( .A(n1414), .B(n1413), .Y(n1419) );
  NOR2XL U1911 ( .A(work_cntr[11]), .B(n1418), .Y(n1412) );
  NAND2XL U1912 ( .A(n1407), .B(n1406), .Y(n1414) );
  NAND2XL U1913 ( .A(n1411), .B(n215), .Y(n1406) );
  NAND2BXL U1914 ( .AN(n1407), .B(n1408), .Y(n1413) );
  NAND2XL U1915 ( .A(n1403), .B(n1405), .Y(n1408) );
  NAND2XL U1916 ( .A(n1402), .B(n1401), .Y(n1405) );
  NAND2XL U1917 ( .A(n1400), .B(n1404), .Y(n1399) );
  NOR2XL U1918 ( .A(work_cntr[13]), .B(n1400), .Y(n1398) );
  NAND2BXL U1919 ( .AN(n1391), .B(n1394), .Y(n1393) );
  INVXL U1920 ( .A(n1387), .Y(n1389) );
  NAND2XL U1921 ( .A(n1386), .B(n1391), .Y(n1392) );
  NAND3XL U1922 ( .A(n1385), .B(n1387), .C(n181), .Y(n1383) );
  NOR2XL U1923 ( .A(work_cntr[15]), .B(n1382), .Y(n1384) );
  NAND2XL U1924 ( .A(n1397), .B(n219), .Y(n1386) );
  AND2XL U1925 ( .A(n1385), .B(n181), .Y(n1379) );
  NAND2XL U1926 ( .A(n182), .B(n128), .Y(n1376) );
  OAI31XL U1927 ( .A0(n1375), .A1(n1381), .A2(n177), .B0(n1380), .Y(n1378) );
  INVXL U1928 ( .A(n1784), .Y(n1380) );
  NOR4X1 U1929 ( .A(write_cntr[13]), .B(write_cntr[12]), .C(write_cntr[14]), 
        .D(n749), .Y(n750) );
  NAND2XL U1930 ( .A(write_cntr[14]), .B(n1522), .Y(n1518) );
  NAND4XL U1931 ( .A(n1756), .B(n1755), .C(n234), .D(n1754), .Y(n1758) );
  AND2XL U1932 ( .A(n2112), .B(n234), .Y(n327) );
  NAND2XL U1933 ( .A(n1506), .B(n234), .Y(n1509) );
  CLKBUFX3 U1934 ( .A(n2347), .Y(en_fb_addr) );
  NAND4BBXL U1935 ( .AN(global_cntr[18]), .BN(global_cntr[5]), .C(n1512), .D(
        n255), .Y(n1513) );
  NOR4XL U1936 ( .A(global_cntr[17]), .B(global_cntr[16]), .C(global_cntr[14]), 
        .D(global_cntr[9]), .Y(n1512) );
  MX2XL U1937 ( .A(n2319), .B(n2320), .S0(curr_photo[0]), .Y(next_photo[0]) );
  AOI221XL U1938 ( .A0(n240), .A1(photo_num[1]), .B0(photo_num[0]), .B1(n188), 
        .C0(n2317), .Y(n2318) );
  OAI21XL U1939 ( .A0(cr_read_cntr[3]), .A1(n500), .B0(n501), .Y(N32) );
  OAI22XL U1940 ( .A0(n360), .A1(n2339), .B0(n2338), .B1(n233), .Y(n518) );
  AOI211XL U1941 ( .A0(n2330), .A1(n2329), .B0(n167), .C0(n234), .Y(n2332) );
  OAI21XL U1942 ( .A0(n273), .A1(n108), .B0(n333), .Y(n475) );
  OAI21XL U1943 ( .A0(n273), .A1(n582), .B0(n357), .Y(n473) );
  OAI21XL U1944 ( .A0(n594), .A1(n273), .B0(n336), .Y(n476) );
  OAI21XL U1945 ( .A0(n273), .A1(n586), .B0(n356), .Y(n474) );
  OAI2BB2XL U1946 ( .B0(n273), .B1(n1771), .A0N(n273), .A1N(write_cntr[4]), 
        .Y(n535) );
  OAI21XL U1947 ( .A0(n682), .A1(n259), .B0(n363), .Y(n498) );
  OAI211XL U1948 ( .A0(N1232), .A1(N1233), .B0(n2292), .C0(n2302), .Y(n363) );
  AOI221XL U1949 ( .A0(n256), .A1(n189), .B0(n2296), .B1(n189), .C0(n2298), 
        .Y(n494) );
  OAI21XL U1950 ( .A0(n686), .A1(n654), .B0(n359), .Y(n490) );
  OAI22XL U1951 ( .A0(n2306), .A1(n258), .B0(n2305), .B1(n2304), .Y(n491) );
  OAI21XL U1952 ( .A0(n273), .A1(n640), .B0(n338), .Y(n489) );
  OAI21XL U1953 ( .A0(n273), .A1(n2308), .B0(n339), .Y(n487) );
  OAI21XL U1954 ( .A0(n273), .A1(n2309), .B0(n340), .Y(n486) );
  OAI21XL U1955 ( .A0(n273), .A1(n2311), .B0(n341), .Y(n485) );
  OAI21XL U1956 ( .A0(n273), .A1(n2312), .B0(n342), .Y(n484) );
  OAI21XL U1957 ( .A0(n273), .A1(n615), .B0(n344), .Y(n482) );
  OAI21XL U1958 ( .A0(n600), .A1(n273), .B0(n351), .Y(n478) );
  OAI21XL U1959 ( .A0(n273), .A1(n596), .B0(n353), .Y(n477) );
  CLKINVX1 U1960 ( .A(n2348), .Y(sftr_n[1]) );
  OA22X1 U1961 ( .A0(n1355), .A1(n1341), .B0(n1353), .B1(n1340), .Y(n2307) );
  OA21XL U1962 ( .A0(\intadd_3/SUM[1] ), .A1(n1353), .B0(n1349), .Y(n2309) );
  AOI2BB1X1 U1963 ( .A0N(\intadd_3/SUM[5] ), .A1N(n1353), .B0(n1246), .Y(n615)
         );
  CLKBUFX3 U1964 ( .A(n884), .Y(n270) );
  NOR2X1 U1965 ( .A(next_state[2]), .B(next_state[1]), .Y(n2281) );
  AOI211X1 U1966 ( .A0(n691), .A1(n1764), .B0(n741), .C0(n740), .Y(n743) );
  OAI22XL U1967 ( .A0(n742), .A1(n739), .B0(n276), .B1(n745), .Y(n740) );
  OAI21XL U1968 ( .A0(n203), .A1(n719), .B0(n107), .Y(n720) );
  NOR2X1 U1969 ( .A(n731), .B(n730), .Y(n701) );
  AOI2BB1X1 U1970 ( .A0N(global_cntr[18]), .A1N(n297), .B0(n727), .Y(n692) );
  OR2X1 U1971 ( .A(n288), .B(n195), .Y(n290) );
  XOR2X1 U1972 ( .A(n284), .B(global_cntr[8]), .Y(n702) );
  OA21XL U1973 ( .A0(global_cntr[6]), .A1(n282), .B0(n283), .Y(n704) );
  NOR3X1 U1974 ( .A(n725), .B(n1514), .C(n724), .Y(n726) );
  NAND4XL U1975 ( .A(global_cntr[19]), .B(global_cntr[16]), .C(global_cntr[14]), .D(global_cntr[9]), .Y(n724) );
  NOR4XL U1976 ( .A(global_cntr[6]), .B(global_cntr[7]), .C(global_cntr[8]), 
        .D(global_cntr[10]), .Y(n722) );
  NOR4XL U1977 ( .A(global_cntr[11]), .B(global_cntr[12]), .C(global_cntr[13]), 
        .D(global_cntr[15]), .Y(n723) );
  NAND2XL U1978 ( .A(global_cntr[18]), .B(global_cntr[17]), .Y(n725) );
  OA21XL U1979 ( .A0(global_cntr[10]), .A1(n287), .B0(n288), .Y(n700) );
  OR2X1 U1980 ( .A(n286), .B(n197), .Y(n288) );
  CLKBUFX3 U1981 ( .A(N582), .Y(n272) );
  AOI21X1 U1982 ( .A0(n669), .A1(n664), .B0(n331), .Y(n662) );
  NOR2X1 U1983 ( .A(n329), .B(n716), .Y(n2348) );
  AOI2BB1X1 U1984 ( .A0N(n1506), .A1N(n234), .B0(n1505), .Y(n1507) );
  OAI21XL U1985 ( .A0(n1504), .A1(n1503), .B0(n1502), .Y(n1505) );
  OA21XL U1986 ( .A0(n187), .A1(n1501), .B0(n1497), .Y(n1506) );
  OAI22XL U1987 ( .A0(n2314), .A1(n232), .B0(im_wen_n), .B1(n574), .Y(n471) );
  OAI22XL U1988 ( .A0(n2314), .A1(n252), .B0(n2313), .B1(im_wen_n), .Y(n472)
         );
  OA21XL U1989 ( .A0(cr_read_cntr[3]), .A1(n2294), .B0(n2295), .Y(n496) );
  OAI21XL U1990 ( .A0(n241), .A1(n2314), .B0(n343), .Y(n483) );
  OAI21XL U1991 ( .A0(n2314), .A1(n243), .B0(n346), .Y(n480) );
  OAI21XL U1992 ( .A0(n245), .A1(n2314), .B0(n350), .Y(n479) );
  CLKINVX1 U1993 ( .A(n1353), .Y(n689) );
  NOR2BX1 U1994 ( .AN(n2278), .B(n14), .Y(n299) );
  AO21X1 U1995 ( .A0(state[0]), .A1(n2316), .B0(n742), .Y(n737) );
  NAND2X1 U1996 ( .A(n291), .B(global_cntr[13]), .Y(n293) );
  NAND2X1 U1997 ( .A(n691), .B(n367), .Y(n329) );
  AO22X1 U1998 ( .A0(n2319), .A1(n366), .B0(curr_photo[1]), .B1(n2320), .Y(
        next_photo[1]) );
  OAI2BB1X1 U1999 ( .A0N(n928), .A1N(n431), .B0(n430), .Y(n432) );
  AO22X1 U2000 ( .A0(n462), .A1(n424), .B0(n461), .B1(n423), .Y(n425) );
  OAI22XL U2001 ( .A0(n437), .A1(n422), .B0(n421), .B1(n420), .Y(n424) );
  OAI21XL U2002 ( .A0(n416), .A1(n415), .B0(n414), .Y(n427) );
  OAI21XL U2003 ( .A0(curr_time[9]), .A1(n457), .B0(n413), .Y(n414) );
  OAI22XL U2004 ( .A0(n441), .A1(n440), .B0(n439), .B1(n450), .Y(n442) );
  OAI2BB2XL U2005 ( .B0(n451), .B1(n450), .A0N(n462), .A1N(\s_0[0] ), .Y(n452)
         );
  OAI2BB1X1 U2006 ( .A0N(n398), .A1N(n438), .B0(n420), .Y(n419) );
  OR2X1 U2007 ( .A(n391), .B(n390), .Y(n400) );
  OAI21XL U2008 ( .A0(n925), .A1(n711), .B0(n405), .Y(n407) );
  OAI2BB1X1 U2009 ( .A0N(n312), .A1N(n311), .B0(n310), .Y(n410) );
  AOI2BB2X1 U2010 ( .B0(n309), .B1(n308), .A0N(n923), .A1N(n924), .Y(n313) );
  AOI2BB2X1 U2011 ( .B0(n376), .B1(n378), .A0N(n937), .A1N(n377), .Y(n382) );
  OAI2BB1X1 U2012 ( .A0N(n937), .A1N(n379), .B0(n377), .Y(n435) );
  OAI2BB1X1 U2013 ( .A0N(n375), .A1N(n374), .B0(n373), .Y(n377) );
  OA21XL U2014 ( .A0(n503), .A1(n502), .B0(n501), .Y(N31) );
  NAND3BX1 U2015 ( .AN(n976), .B(n468), .C(n256), .Y(n469) );
  NAND2XL U2016 ( .A(n234), .B(n1608), .Y(n1607) );
  AO21X1 U2017 ( .A0(N1234), .A1(n365), .B0(n364), .Y(n497) );
  NAND3XL U2018 ( .A(n2106), .B(N2062), .C(n187), .Y(n2104) );
  OAI211XL U2019 ( .A0(n2106), .A1(n187), .B0(n2107), .C0(n167), .Y(n2105) );
  OAI2BB1X1 U2020 ( .A0N(n676), .A1N(\C162/DATA3_1 ), .B0(n670), .Y(n671) );
  AOI2BB2X1 U2021 ( .B0(n269), .B1(N1447), .A0N(n254), .A1N(n204), .Y(n670) );
  OAI2BB1X1 U2022 ( .A0N(n676), .A1N(\C162/DATA3_2 ), .B0(n672), .Y(n673) );
  AOI2BB2X1 U2023 ( .B0(n269), .B1(N1448), .A0N(n254), .A1N(n161), .Y(n672) );
  OAI2BB1X1 U2024 ( .A0N(n676), .A1N(\C162/DATA3_17 ), .B0(n674), .Y(n675) );
  AOI2BB2X1 U2025 ( .B0(n269), .B1(N1463), .A0N(n254), .A1N(n202), .Y(n674) );
  OA21XL U2026 ( .A0(n669), .A1(n668), .B0(n223), .Y(n169) );
  OAI22XL U2027 ( .A0(n577), .A1(n660), .B0(n276), .B1(n255), .Y(
        \U3/RSOP_657/C2/Z_19 ) );
  OAI22XL U2028 ( .A0(n578), .A1(n232), .B0(n641), .B1(n574), .Y(n575) );
  OAI22XL U2029 ( .A0(n653), .A1(n660), .B0(n276), .B1(n204), .Y(
        \U3/RSOP_657/C2/Z_1 ) );
  OAI22XL U2030 ( .A0(n649), .A1(n237), .B0(n648), .B1(n238), .Y(n650) );
  OAI2BB2XL U2031 ( .B0(n188), .B1(n276), .A0N(curr_photo_addr[1]), .A1N(n661), 
        .Y(n678) );
  OAI22XL U2032 ( .A0(n659), .A1(n660), .B0(n276), .B1(n236), .Y(
        \U3/RSOP_657/C2/Z_0 ) );
  AOI222XL U2033 ( .A0(n658), .A1(n657), .B0(n656), .B1(\next_write_addr_w[0] ), .C0(n124), .C1(n655), .Y(n659) );
  OAI2BB2XL U2034 ( .B0(n240), .B1(n276), .A0N(curr_photo_addr[2]), .A1N(n661), 
        .Y(n679) );
  OAI22XL U2035 ( .A0(n646), .A1(n660), .B0(n276), .B1(n161), .Y(
        \U3/RSOP_657/C2/Z_2 ) );
  OAI22XL U2036 ( .A0(n649), .A1(n238), .B0(n648), .B1(n235), .Y(n643) );
  OAI2BB1X1 U2037 ( .A0N(curr_photo_addr[3]), .A1N(n661), .B0(n2334), .Y(n680)
         );
  OAI22XL U2038 ( .A0(n639), .A1(n660), .B0(n276), .B1(n242), .Y(
        \U3/RSOP_657/C2/Z_3 ) );
  OAI22XL U2039 ( .A0(n649), .A1(n235), .B0(n648), .B1(n162), .Y(n636) );
  OA21XL U2040 ( .A0(n265), .A1(n235), .B0(n2307), .Y(n642) );
  OAI2BB1X1 U2041 ( .A0N(curr_photo_addr[4]), .A1N(n661), .B0(n2334), .Y(
        \C1/Z_4 ) );
  OAI22XL U2042 ( .A0(n635), .A1(n660), .B0(n276), .B1(n190), .Y(
        \U3/RSOP_657/C2/Z_4 ) );
  OAI22XL U2043 ( .A0(n649), .A1(n162), .B0(n648), .B1(n239), .Y(n633) );
  OAI22XL U2044 ( .A0(n631), .A1(n660), .B0(n276), .B1(n630), .Y(
        \U3/RSOP_657/C2/Z_5 ) );
  OAI22XL U2045 ( .A0(n649), .A1(n239), .B0(n648), .B1(n2310), .Y(n627) );
  OA21XL U2046 ( .A0(n265), .A1(n239), .B0(n2309), .Y(n632) );
  OAI22XL U2047 ( .A0(n626), .A1(n660), .B0(n276), .B1(n196), .Y(
        \U3/RSOP_657/C2/Z_6 ) );
  OAI22XL U2048 ( .A0(n649), .A1(n2310), .B0(n648), .B1(n163), .Y(n624) );
  OAI2BB1X1 U2049 ( .A0N(curr_photo_addr[7]), .A1N(n661), .B0(n2334), .Y(
        \C1/Z_7 ) );
  OAI22XL U2050 ( .A0(n622), .A1(n660), .B0(n276), .B1(n194), .Y(
        \U3/RSOP_657/C2/Z_7 ) );
  OAI22XL U2051 ( .A0(n649), .A1(n163), .B0(n648), .B1(n241), .Y(n619) );
  OA21XL U2052 ( .A0(n265), .A1(n163), .B0(n2312), .Y(n623) );
  OAI22XL U2053 ( .A0(n618), .A1(n660), .B0(n276), .B1(n200), .Y(
        \U3/RSOP_657/C2/Z_8 ) );
  OAI22XL U2054 ( .A0(n649), .A1(n241), .B0(n648), .B1(n165), .Y(n616) );
  AO22X1 U2055 ( .A0(n614), .A1(n613), .B0(n171), .B1(global_cntr[9]), .Y(
        \U3/RSOP_657/C2/Z_9 ) );
  OAI222XL U2056 ( .A0(n244), .A1(n648), .B0(n641), .B1(n612), .C0(n2330), 
        .C1(n233), .Y(n613) );
  OAI22XL U2057 ( .A0(n611), .A1(n660), .B0(n276), .B1(n197), .Y(
        \U3/RSOP_657/C2/Z_10 ) );
  OAI22XL U2058 ( .A0(n649), .A1(n165), .B0(n648), .B1(n243), .Y(n608) );
  OAI2BB1X1 U2059 ( .A0N(curr_photo_addr[11]), .A1N(n661), .B0(n2334), .Y(
        \C1/Z_11 ) );
  OAI22XL U2060 ( .A0(n607), .A1(n660), .B0(n276), .B1(n195), .Y(
        \U3/RSOP_657/C2/Z_11 ) );
  OAI22XL U2061 ( .A0(n649), .A1(n244), .B0(n648), .B1(n245), .Y(n604) );
  OAI22XL U2062 ( .A0(n603), .A1(n660), .B0(n276), .B1(n198), .Y(
        \U3/RSOP_657/C2/Z_12 ) );
  OAI22XL U2063 ( .A0(n649), .A1(n243), .B0(n164), .B1(n648), .Y(n601) );
  AOI2BB1X1 U2064 ( .A0N(n1243), .A1N(n1355), .B0(n1244), .Y(n345) );
  OAI2BB1X1 U2065 ( .A0N(curr_photo_addr[13]), .A1N(n661), .B0(n2334), .Y(
        \C1/Z_13 ) );
  OAI22XL U2066 ( .A0(n599), .A1(n660), .B0(n276), .B1(n250), .Y(
        \U3/RSOP_657/C2/Z_13 ) );
  OAI22XL U2067 ( .A0(n649), .A1(n245), .B0(n648), .B1(n166), .Y(n597) );
  OAI2BB1X1 U2068 ( .A0N(n689), .A1N(\intadd_4/SUM[2] ), .B0(n349), .Y(n606)
         );
  OAI2BB1X1 U2069 ( .A0N(curr_photo_addr[14]), .A1N(n661), .B0(n2334), .Y(
        \C1/Z_14 ) );
  OAI2BB1X1 U2070 ( .A0N(curr_photo_addr[15]), .A1N(n661), .B0(n2334), .Y(
        \C1/Z_15 ) );
  OAI22XL U2071 ( .A0(n593), .A1(n660), .B0(n276), .B1(n199), .Y(
        \U3/RSOP_657/C2/Z_15 ) );
  OAI22XL U2072 ( .A0(n108), .A1(n641), .B0(n648), .B1(n247), .Y(n590) );
  OAI22XL U2073 ( .A0(n589), .A1(n660), .B0(n276), .B1(n251), .Y(
        \U3/RSOP_657/C2/Z_16 ) );
  OAI22XL U2074 ( .A0(n586), .A1(n641), .B0(n648), .B1(n248), .Y(n587) );
  AO21X1 U2075 ( .A0(n718), .A1(n334), .B0(n1313), .Y(n335) );
  OAI22XL U2076 ( .A0(n585), .A1(n660), .B0(n276), .B1(n202), .Y(
        \U3/RSOP_657/C2/Z_17 ) );
  OAI22XL U2077 ( .A0(n582), .A1(n641), .B0(n648), .B1(n231), .Y(n583) );
  OAI2BB1X1 U2078 ( .A0N(n1371), .A1N(n1362), .B0(n512), .Y(n513) );
  AOI2BB2X1 U2079 ( .B0(n511), .B1(n1370), .A0N(n1362), .A1N(n510), .Y(n514)
         );
  OR2X1 U2080 ( .A(n1308), .B(n358), .Y(n574) );
  OAI22XL U2081 ( .A0(n1333), .A1(n232), .B0(n1335), .B1(n1334), .Y(n358) );
  OAI22XL U2082 ( .A0(n581), .A1(n660), .B0(n276), .B1(n253), .Y(
        \U3/RSOP_657/C2/Z_18 ) );
  OAI22XL U2083 ( .A0(n578), .A1(n252), .B0(n2313), .B1(n641), .Y(n579) );
  AOI2BB1X1 U2084 ( .A0N(n265), .A1N(n641), .B0(n656), .Y(n578) );
  OA21XL U2085 ( .A0(global_cntr[11]), .A1(n289), .B0(n290), .Y(n699) );
  OA21XL U2086 ( .A0(global_cntr[3]), .A1(n708), .B0(n280), .Y(n707) );
  OA21XL U2087 ( .A0(global_cntr[5]), .A1(n281), .B0(n729), .Y(n705) );
  OA21XL U2088 ( .A0(global_cntr[13]), .A1(n291), .B0(n293), .Y(n697) );
  OAI2BB1X1 U2089 ( .A0N(n1195), .A1N(n1510), .B0(n361), .Y(n1368) );
  NAND2XL U2090 ( .A(n2326), .B(n234), .Y(n1195) );
  OAI22XL U2091 ( .A0(n509), .A1(n1370), .B0(n1371), .B1(n233), .Y(n566) );
  OAI21XL U2092 ( .A0(n1373), .A1(n1605), .B0(n507), .Y(n508) );
  NAND4XL U2093 ( .A(write_addr[9]), .B(write_addr[10]), .C(write_addr[11]), 
        .D(write_addr[12]), .Y(n1357) );
  OAI2BB1X1 U2094 ( .A0N(n665), .A1N(n2348), .B0(n330), .Y(n331) );
  OR2X1 U2095 ( .A(state[0]), .B(n716), .Y(n369) );
  AOI2BB2X1 U2096 ( .B0(n2112), .B1(n326), .A0N(n1373), .A1N(n1374), .Y(n665)
         );
  OA21XL U2097 ( .A0(n885), .A1(n229), .B0(n752), .Y(n174) );
  OA22X1 U2098 ( .A0(n265), .A1(n241), .B0(n1355), .B1(n1354), .Y(n186) );
  OR2X1 U2099 ( .A(n1247), .B(n769), .Y(n193) );
  OA22X1 U2100 ( .A0(n667), .A1(n666), .B0(n665), .B1(sftr_n[1]), .Y(n223) );
  CLKBUFX3 U2101 ( .A(write_addr[17]), .Y(n271) );
  OAI31XL U2102 ( .A0(write_cntr[7]), .A1(write_cntr[5]), .A2(write_cntr[6]), 
        .B0(write_cntr[8]), .Y(n719) );
  OAI31XL U2103 ( .A0(write_cntr[9]), .A1(write_cntr[10]), .A2(n747), .B0(
        write_cntr[11]), .Y(n748) );
  AND4X1 U2104 ( .A(write_cntr[7]), .B(write_cntr[6]), .C(write_cntr[8]), .D(
        n780), .Y(n766) );
  OAI21XL U2105 ( .A0(write_cntr[14]), .A1(n753), .B0(n783), .Y(n752) );
  AOI2BB2X1 U2106 ( .B0(write_cntr[12]), .B1(n755), .A0N(write_cntr[12]), 
        .A1N(n755), .Y(n754) );
  AOI2BB2X1 U2107 ( .B0(n117), .B1(n175), .A0N(n117), .A1N(n175), .Y(n960) );
  AOI221XL U2108 ( .A0(n1777), .A1(n173), .B0(n779), .B1(n173), .C0(n766), .Y(
        n767) );
  AO21X1 U2109 ( .A0(n881), .A1(n208), .B0(n270), .Y(n774) );
  AOI2BB2X1 U2110 ( .B0(n1249), .B1(n964), .A0N(n1249), .A1N(n964), .Y(n806)
         );
  AOI2BB2X1 U2111 ( .B0(n794), .B1(n793), .A0N(n794), .A1N(n793), .Y(n807) );
  OAI21XL U2112 ( .A0(n799), .A1(n796), .B0(n798), .Y(n797) );
  OAI21XL U2113 ( .A0(n819), .A1(n823), .B0(n818), .Y(n817) );
  AOI2BB2X1 U2114 ( .B0(n1256), .B1(n115), .A0N(n1256), .A1N(n115), .Y(n828)
         );
  AOI2BB2X1 U2115 ( .B0(n1778), .B1(n1264), .A0N(n1778), .A1N(n1264), .Y(n841)
         );
  OR2X1 U2116 ( .A(n841), .B(n1023), .Y(n845) );
  OAI21XL U2117 ( .A0(n834), .A1(n1264), .B0(n833), .Y(n831) );
  AOI2BB2X1 U2118 ( .B0(n1023), .B1(n1268), .A0N(n1023), .A1N(n1268), .Y(n851)
         );
  OAI31XL U2119 ( .A0(n842), .A1(n1023), .A2(n841), .B0(n840), .Y(n843) );
  AOI2BB2X1 U2120 ( .B0(n1277), .B1(n1775), .A0N(n1277), .A1N(n1775), .Y(n865)
         );
  OAI2BB1X1 U2121 ( .A0N(n855), .A1N(n854), .B0(n857), .Y(n856) );
  AOI2BB2X1 U2122 ( .B0(n1771), .B1(n1280), .A0N(n1771), .A1N(n1280), .Y(n887)
         );
  OAI2BB1X1 U2123 ( .A0N(n868), .A1N(n867), .B0(n870), .Y(n869) );
  OAI2BB1X1 U2124 ( .A0N(n877), .A1N(n886), .B0(n879), .Y(n878) );
  OAI21XL U2125 ( .A0(n882), .A1(write_cntr[2]), .B0(n881), .Y(n883) );
  AOI2BB2X1 U2126 ( .B0(n1301), .B1(n1774), .A0N(n1301), .A1N(n1774), .Y(n900)
         );
  OAI21XL U2127 ( .A0(n1288), .A1(n895), .B0(n896), .Y(n894) );
  OAI21XL U2128 ( .A0(n905), .A1(n1288), .B0(n904), .Y(n902) );
  OAI31XL U2129 ( .A0(n905), .A1(n904), .A2(n903), .B0(n902), .Y(n906) );
  OR2X1 U2130 ( .A(n915), .B(n916), .Y(n907) );
  AOI2BB2X1 U2131 ( .B0(n1769), .B1(n1240), .A0N(n1769), .A1N(n1240), .Y(n1199) );
  AOI2BB2X1 U2132 ( .B0(n909), .B1(n908), .A0N(n909), .A1N(n908), .Y(n1205) );
  OAI21XL U2133 ( .A0(n913), .A1(n1240), .B0(n912), .Y(n910) );
  OAI21XL U2134 ( .A0(n1240), .A1(n915), .B0(n916), .Y(n914) );
  AOI2BB1X1 U2135 ( .A0N(work_cntr[10]), .A1N(n949), .B0(n950), .Y(n1851) );
  AOI2BB2X1 U2136 ( .B0(n215), .B1(n951), .A0N(n215), .A1N(n951), .Y(n1829) );
  AOI2BB1X1 U2137 ( .A0N(work_cntr[15]), .A1N(n954), .B0(n955), .Y(n1798) );
  AO21X1 U2138 ( .A0(n213), .A1(n1783), .B0(n956), .Y(n1959) );
  AOI2BB2X1 U2139 ( .B0(work_cntr[19]), .B1(n1785), .A0N(work_cntr[19]), .A1N(
        n1785), .Y(n1967) );
  NAND3BX1 U2140 ( .AN(n998), .B(n1002), .C(n1010), .Y(n999) );
  AOI2BB2X1 U2141 ( .B0(n232), .B1(n1055), .A0N(n232), .A1N(n1055), .Y(n1334)
         );
  AO21X1 U2142 ( .A0(n983), .A1(n164), .B0(n984), .Y(n1304) );
  AOI2BB2X1 U2143 ( .B0(n1336), .B1(n162), .A0N(n1336), .A1N(n162), .Y(n1346)
         );
  AOI2BB2X1 U2144 ( .B0(n1347), .B1(n2310), .A0N(n1347), .A1N(n2310), .Y(n1350) );
  AOI2BB2X1 U2145 ( .B0(n987), .B1(N584), .A0N(n987), .A1N(N584), .Y(n1351) );
  AOI2BB2X1 U2146 ( .B0(n1001), .B1(n1000), .A0N(n1001), .A1N(n1000), .Y(n1015) );
  AOI2BB2X1 U2147 ( .B0(n1012), .B1(n1007), .A0N(n1012), .A1N(n1007), .Y(n1022) );
  AO22X1 U2148 ( .A0(n1778), .A1(n1217), .B0(n1008), .B1(n1024), .Y(n1009) );
  AOI2BB2X1 U2149 ( .B0(n1024), .B1(n1036), .A0N(n1023), .A1N(n1231), .Y(n1025) );
  AOI2BB2X1 U2150 ( .B0(n1026), .B1(n1025), .A0N(n1026), .A1N(n1025), .Y(n1046) );
  AOI2BB2X1 U2151 ( .B0(n1030), .B1(n1029), .A0N(n1030), .A1N(n1029), .Y(n1052) );
  AOI2BB2X1 U2152 ( .B0(n1039), .B1(n1038), .A0N(n1039), .A1N(n1038), .Y(n1044) );
  OAI21XL U2153 ( .A0(\intadd_3/A[0] ), .A1(n1771), .B0(n1040), .Y(n1041) );
  OAI22XL U2154 ( .A0(n1046), .A1(n1047), .B0(n1044), .B1(n1043), .Y(n1045) );
  OAI2BB1X1 U2155 ( .A0N(n1047), .A1N(n1046), .B0(n1045), .Y(n1053) );
  AOI2BB2X1 U2156 ( .B0(n1065), .B1(n1297), .A0N(n1065), .A1N(n1297), .Y(n1057) );
  AOI2BB2X1 U2157 ( .B0(n1058), .B1(\next_write_addr_w[0] ), .A0N(n1058), 
        .A1N(n1057), .Y(n1062) );
  OAI21XL U2158 ( .A0(n1060), .A1(n1059), .B0(n1297), .Y(n1061) );
  OAI22XL U2159 ( .A0(n1355), .A1(n1062), .B0(n1327), .B1(n1061), .Y(n1063) );
  NOR2X1 U2160 ( .A(work_cntr[19]), .B(n1068), .Y(n2321) );
  AO21X1 U2161 ( .A0(n1075), .A1(work_cntr[16]), .B0(n1066), .Y(n1081) );
  AOI2BB2X1 U2162 ( .B0(n1081), .B1(n1080), .A0N(n1081), .A1N(n1080), .Y(n1085) );
  OAI2BB1X1 U2163 ( .A0N(work_cntr[16]), .A1N(n1080), .B0(n1079), .Y(n1090) );
  OR2X1 U2164 ( .A(n1081), .B(n1080), .Y(n1083) );
  AO21X1 U2165 ( .A0(n181), .A1(n1094), .B0(n1086), .Y(n1084) );
  AOI2BB2X1 U2166 ( .B0(n1085), .B1(n1091), .A0N(n1085), .A1N(n1084), .Y(n1092) );
  OAI2BB1X1 U2167 ( .A0N(n1091), .A1N(n1090), .B0(n1089), .Y(n1093) );
  OR2X1 U2168 ( .A(n1093), .B(n1092), .Y(n1105) );
  OAI21XL U2169 ( .A0(work_cntr[13]), .A1(n1108), .B0(n1099), .Y(n1097) );
  AOI2BB2X1 U2170 ( .B0(work_cntr[13]), .B1(n1096), .A0N(work_cntr[13]), .A1N(
        n1096), .Y(n1107) );
  NAND3BX1 U2171 ( .AN(n1115), .B(n1101), .C(n1108), .Y(n1100) );
  AO21X1 U2172 ( .A0(work_cntr[11]), .A1(n1103), .B0(n1102), .Y(n1121) );
  OAI21XL U2173 ( .A0(n1105), .A1(n219), .B0(n1104), .Y(n1106) );
  OAI21XL U2174 ( .A0(work_cntr[12]), .A1(n1121), .B0(n1114), .Y(n1109) );
  AO21X1 U2175 ( .A0(n222), .A1(n1123), .B0(n1122), .Y(n1111) );
  OA22X1 U2176 ( .A0(n1113), .A1(n1121), .B0(n1112), .B1(n1111), .Y(n1119) );
  NAND3BX1 U2177 ( .AN(n1117), .B(n1121), .C(n1122), .Y(n1120) );
  OAI21XL U2178 ( .A0(work_cntr[9]), .A1(n1133), .B0(n1131), .Y(n1129) );
  NAND3BX1 U2179 ( .AN(n1146), .B(n1134), .C(n1133), .Y(n1132) );
  AO21X1 U2180 ( .A0(work_cntr[7]), .A1(n1136), .B0(n1135), .Y(n1155) );
  OAI2BB1X1 U2181 ( .A0N(n1156), .A1N(work_cntr[6]), .B0(n1136), .Y(n1159) );
  OAI21XL U2182 ( .A0(n183), .A1(n1138), .B0(n1137), .Y(n1139) );
  OAI21XL U2183 ( .A0(work_cntr[8]), .A1(n1155), .B0(n1148), .Y(n1141) );
  OAI21XL U2184 ( .A0(work_cntr[7]), .A1(n1159), .B0(n1154), .Y(n1143) );
  NOR3BXL U2185 ( .AN(n1155), .B(n1152), .C(n1154), .Y(n1149) );
  NAND3BX1 U2186 ( .AN(n1149), .B(n1151), .C(n1159), .Y(n1150) );
  OAI21XL U2187 ( .A0(n1152), .A1(n1154), .B0(n1155), .Y(n1153) );
  OAI21XL U2188 ( .A0(work_cntr[6]), .A1(n1171), .B0(n1158), .Y(n1161) );
  OAI31XL U2189 ( .A0(n1177), .A1(work_cntr[5]), .A2(n1166), .B0(n1165), .Y(
        n1167) );
  OA21XL U2190 ( .A0(n1175), .A1(n1174), .B0(n1177), .Y(n1176) );
  AOI2BB2X1 U2191 ( .B0(n1178), .B1(n1177), .A0N(n1178), .A1N(n1176), .Y(n1183) );
  OAI21XL U2192 ( .A0(n1922), .A1(n1911), .B0(n1183), .Y(n1179) );
  AOI2BB2X1 U2193 ( .B0(n1922), .B1(n109), .A0N(n1922), .A1N(n109), .Y(n1190)
         );
  OAI21XL U2194 ( .A0(n1181), .A1(n1183), .B0(n1911), .Y(n1182) );
  OAI2BB1X1 U2195 ( .A0N(n1934), .A1N(n109), .B0(n1922), .Y(n1187) );
  OAI21XL U2196 ( .A0(n1194), .A1(n1191), .B0(n1939), .Y(n1189) );
  AOI2BB2X1 U2197 ( .B0(n1190), .B1(n1189), .A0N(n1190), .A1N(n1934), .Y(n2327) );
  AOI2BB2X1 U2198 ( .B0(n114), .B1(n1209), .A0N(n114), .A1N(n1209), .Y(n1201)
         );
  AOI222XL U2199 ( .A0(\intadd_3/B[0] ), .A1(n132), .B0(\intadd_3/B[0] ), .B1(
        n131), .C0(n132), .C1(n131), .Y(n1343) );
  AOI2BB1X1 U2200 ( .A0N(n1218), .A1N(n1237), .B0(n1227), .Y(n1220) );
  ADDFXL U2201 ( .A(n1224), .B(n1221), .CI(n1220), .CO(n1222), .S(n1219) );
  AOI2BB1X1 U2202 ( .A0N(n1224), .A1N(next_cr_x[5]), .B0(n1234), .Y(n1226) );
  ADDFXL U2203 ( .A(n1231), .B(n1227), .CI(n1226), .CO(n1228), .S(n1225) );
  AOI2BB1X1 U2204 ( .A0N(n1231), .A1N(next_cr_x[6]), .B0(n1238), .Y(n1233) );
  ADDFXL U2205 ( .A(n1237), .B(n1234), .CI(n1233), .CO(n1235), .S(n1232) );
  ADDFXL U2206 ( .A(next_cr_x[5]), .B(n1238), .CI(n1237), .CO(n1239), .S(n1236) );
  OAI2BB1X1 U2207 ( .A0N(n1247), .A1N(n1248), .B0(n1248), .Y(n1254) );
  AOI2BB2X1 U2208 ( .B0(n1257), .B1(n1255), .A0N(n1257), .A1N(n1255), .Y(n1263) );
  AOI2BB2X1 U2209 ( .B0(n1254), .B1(n1253), .A0N(n1254), .A1N(n1252), .Y(n1259) );
  AOI2BB2X1 U2210 ( .B0(n1259), .B1(n1258), .A0N(n1259), .A1N(n1257), .Y(n1267) );
  OAI21XL U2211 ( .A0(n1261), .A1(n1263), .B0(n1265), .Y(n1262) );
  AOI2BB2X1 U2212 ( .B0(n1276), .B1(n1274), .A0N(n1276), .A1N(n1273), .Y(n1283) );
  AOI2BB2X1 U2213 ( .B0(n1277), .B1(n1275), .A0N(n1277), .A1N(n1275), .Y(n1284) );
  AOI222XL U2214 ( .A0(n1320), .A1(n1319), .B0(n1320), .B1(n718), .C0(n1319), 
        .C1(n1318), .Y(n1321) );
  OAI21XL U2215 ( .A0(N580), .A1(N579), .B0(n1336), .Y(n1341) );
  AOI2BB2X1 U2216 ( .B0(n132), .B1(n131), .A0N(n132), .A1N(n131), .Y(n1339) );
  AOI2BB2X1 U2217 ( .B0(\intadd_3/B[0] ), .B1(n1339), .A0N(\intadd_3/B[0] ), 
        .A1N(n1339), .Y(n1340) );
  ADDFXL U2218 ( .A(n1344), .B(n1343), .CI(n1342), .CO(n1216), .S(n1345) );
  AOI2BB2X1 U2219 ( .B0(n1350), .B1(n718), .A0N(\intadd_3/SUM[2] ), .A1N(n1353), .Y(n2311) );
  AOI2BB2X1 U2220 ( .B0(n1351), .B1(n718), .A0N(\intadd_3/SUM[3] ), .A1N(n1353), .Y(n2312) );
  OAI21XL U2221 ( .A0(n1365), .A1(n1511), .B0(n684), .Y(n1366) );
  AO21X1 U2222 ( .A0(n212), .A1(work_cntr[17]), .B0(n1375), .Y(n1377) );
  AO21X1 U2223 ( .A0(work_cntr[18]), .A1(n1381), .B0(n1784), .Y(n1387) );
  AOI2BB2X1 U2224 ( .B0(work_cntr[15]), .B1(n1382), .A0N(work_cntr[15]), .A1N(
        n1382), .Y(n1397) );
  AO21X1 U2225 ( .A0(n1390), .A1(n1389), .B0(n1388), .Y(n1394) );
  OAI2BB1X1 U2226 ( .A0N(n1392), .A1N(n1394), .B0(n219), .Y(n1396) );
  OAI21XL U2227 ( .A0(n1394), .A1(work_cntr[14]), .B0(n1397), .Y(n1395) );
  OR2X1 U2228 ( .A(n1398), .B(n1402), .Y(n1403) );
  OAI2BB1X1 U2229 ( .A0N(n1403), .A1N(n1401), .B0(n221), .Y(n1404) );
  OA21XL U2230 ( .A0(n221), .A1(n1405), .B0(n1404), .Y(n1411) );
  OAI2BB1X1 U2231 ( .A0N(n1414), .A1N(n1408), .B0(n215), .Y(n1410) );
  OAI21XL U2232 ( .A0(n1408), .A1(work_cntr[12]), .B0(n1411), .Y(n1409) );
  OR2X1 U2233 ( .A(n1412), .B(n122), .Y(n1416) );
  OAI2BB1X1 U2234 ( .A0N(n1416), .A1N(n1419), .B0(n222), .Y(n1421) );
  OAI21XL U2235 ( .A0(n1419), .A1(work_cntr[11]), .B0(n1422), .Y(n1420) );
  OAI2BB1X1 U2236 ( .A0N(n1437), .A1N(n1433), .B0(n214), .Y(n1434) );
  AOI2BB1X1 U2237 ( .A0N(n226), .A1N(n1443), .B0(n1442), .Y(n1452) );
  OAI21XL U2238 ( .A0(n1449), .A1(work_cntr[7]), .B0(n1452), .Y(n1450) );
  OAI2BB1X1 U2239 ( .A0N(n1464), .A1N(n1466), .B0(n168), .Y(n1468) );
  OAI21XL U2240 ( .A0(n1466), .A1(work_cntr[5]), .B0(n1469), .Y(n1467) );
  OR2X1 U2241 ( .A(n1470), .B(n1474), .Y(n1475) );
  OAI2BB1X1 U2242 ( .A0N(n1475), .A1N(n1473), .B0(n180), .Y(n1476) );
  OA21XL U2243 ( .A0(n180), .A1(n1477), .B0(n1476), .Y(n1483) );
  OAI2BB1X1 U2244 ( .A0N(n1487), .A1N(n1480), .B0(n179), .Y(n1482) );
  OAI21XL U2245 ( .A0(n1480), .A1(N2063), .B0(n1483), .Y(n1481) );
  OR2X1 U2246 ( .A(n119), .B(n1485), .Y(n1492) );
  OAI2BB1X1 U2247 ( .A0N(n1492), .A1N(n1490), .B0(n167), .Y(n1493) );
  OAI21XL U2248 ( .A0(n1490), .A1(N2062), .B0(n1489), .Y(n1488) );
  OAI2BB1X1 U2249 ( .A0N(n1500), .A1N(n1499), .B0(n1502), .Y(n1508) );
  NAND3BX1 U2250 ( .AN(write_cntr[12]), .B(n230), .C(n1519), .Y(n1522) );
  AOI2BB2X1 U2251 ( .B0(write_cntr[12]), .B1(n1521), .A0N(write_cntr[12]), 
        .A1N(n1521), .Y(n1530) );
  NAND3BX1 U2252 ( .AN(n130), .B(n1530), .C(n1526), .Y(n1533) );
  AOI2BB2X1 U2253 ( .B0(n130), .B1(n1527), .A0N(n130), .A1N(n1527), .Y(n1544)
         );
  NAND3BX1 U2254 ( .AN(n1542), .B(n1544), .C(n1535), .Y(n1547) );
  OA22X1 U2255 ( .A0(n1534), .A1(n1533), .B0(n1532), .B1(n1531), .Y(n1545) );
  AOI2BB2X1 U2256 ( .B0(n1542), .B1(n1541), .A0N(n1542), .A1N(n1541), .Y(n1551) );
  NAND3BX1 U2257 ( .AN(n1558), .B(n1551), .C(n1549), .Y(n1561) );
  OA22X1 U2258 ( .A0(n1548), .A1(n1547), .B0(n1546), .B1(n1545), .Y(n1559) );
  AOI2BB2X1 U2259 ( .B0(n1558), .B1(n1557), .A0N(n1558), .A1N(n1557), .Y(n1573) );
  NAND3BX1 U2260 ( .AN(n1571), .B(n1573), .C(n1564), .Y(n1576) );
  NAND4BBXL U2261 ( .AN(n1592), .BN(n1566), .C(write_cntr[4]), .D(n1567), .Y(
        n1585) );
  OR2X1 U2262 ( .A(n1567), .B(n1566), .Y(n1568) );
  AOI2BB2X1 U2263 ( .B0(n1577), .B1(n1576), .A0N(n1577), .A1N(n1575), .Y(n1584) );
  OAI21XL U2264 ( .A0(n1584), .A1(n1586), .B0(n1583), .Y(n1600) );
  OAI21XL U2265 ( .A0(write_cntr[4]), .A1(n1767), .B0(write_cntr[3]), .Y(n1589) );
  OAI221XL U2266 ( .A0(n1592), .A1(n1589), .B0(n1593), .B1(n1592), .C0(n1591), 
        .Y(n1590) );
  OAI31XL U2267 ( .A0(n1593), .A1(n1592), .A2(n1591), .B0(n1590), .Y(n1594) );
  OAI2BB1X1 U2268 ( .A0N(n1598), .A1N(n1597), .B0(n1594), .Y(n1595) );
  AO21X1 U2269 ( .A0(work_cntr[11]), .A1(n1611), .B0(n1612), .Y(n1664) );
  AO21X1 U2270 ( .A0(n1615), .A1(n1622), .B0(n1618), .Y(n1616) );
  OAI2BB2XL U2271 ( .B0(n1617), .B1(n1618), .A0N(n1617), .A1N(n1616), .Y(n1625) );
  OR2X1 U2272 ( .A(n1624), .B(n1638), .Y(n1627) );
  AO21X1 U2273 ( .A0(n1625), .A1(n1637), .B0(n1624), .Y(n1630) );
  AO21X1 U2274 ( .A0(n1629), .A1(n1628), .B0(n1627), .Y(n1641) );
  AO21X1 U2275 ( .A0(work_cntr[13]), .A1(n1634), .B0(n1969), .Y(n1645) );
  OAI21XL U2276 ( .A0(n1639), .A1(n1638), .B0(n1637), .Y(n1640) );
  OAI31XL U2277 ( .A0(n1642), .A1(n1641), .A2(n1661), .B0(n1640), .Y(n1644) );
  AOI2BB1X1 U2278 ( .A0N(n1648), .A1N(n1644), .B0(n1643), .Y(n1646) );
  OAI21XL U2279 ( .A0(n1654), .A1(n1655), .B0(n1656), .Y(n1647) );
  OAI21XL U2280 ( .A0(n1661), .A1(n1656), .B0(n1649), .Y(n1650) );
  AOI2BB2X1 U2281 ( .B0(n1654), .B1(n1657), .A0N(n1654), .A1N(n1657), .Y(n1679) );
  OAI21XL U2282 ( .A0(n1662), .A1(n1660), .B0(n1661), .Y(n1659) );
  AOI2BB2X1 U2283 ( .B0(n1666), .B1(n1665), .A0N(n1666), .A1N(n1665), .Y(n1669) );
  NAND3BX1 U2284 ( .AN(n1697), .B(n1686), .C(n1700), .Y(n1691) );
  AOI2BB2X1 U2285 ( .B0(n1688), .B1(n1697), .A0N(n1688), .A1N(n1697), .Y(n1693) );
  OAI21XL U2286 ( .A0(n1700), .A1(n1699), .B0(n1698), .Y(n1703) );
  AOI2BB2X1 U2287 ( .B0(n1707), .B1(n1706), .A0N(n1707), .A1N(n1706), .Y(n1713) );
  AOI221XL U2288 ( .A0(n2122), .A1(n1715), .B0(n1714), .B1(n1715), .C0(n1717), 
        .Y(n1712) );
  OAI2BB1X1 U2289 ( .A0N(n1715), .A1N(n1722), .B0(n1717), .Y(n1716) );
  OR2X1 U2290 ( .A(n1720), .B(n180), .Y(n1726) );
  AOI2BB2X1 U2291 ( .B0(n2122), .B1(n1721), .A0N(n2122), .A1N(n1721), .Y(n1727) );
  AO21X1 U2292 ( .A0(n179), .A1(n1728), .B0(n1727), .Y(n1729) );
  OA22X1 U2293 ( .A0(n1732), .A1(n1731), .B0(n1730), .B1(n1734), .Y(n1743) );
  AOI2BB2X1 U2294 ( .B0(n1752), .B1(n1734), .A0N(n1752), .A1N(n1734), .Y(n1735) );
  OAI22XL U2295 ( .A0(n273), .A1(n1769), .B0(n2314), .B1(n224), .Y(n537) );
  OAI22XL U2296 ( .A0(n273), .A1(n1770), .B0(n2314), .B1(n225), .Y(n536) );
  OAI22XL U2297 ( .A0(n273), .A1(n115), .B0(n2314), .B1(n173), .Y(n534) );
  OAI22XL U2298 ( .A0(n273), .A1(n1773), .B0(n2314), .B1(n185), .Y(n532) );
  OAI22XL U2299 ( .A0(n273), .A1(n1774), .B0(n2314), .B1(n208), .Y(n531) );
  OAI22XL U2300 ( .A0(n273), .A1(n1775), .B0(n2314), .B1(n210), .Y(n530) );
  OAI22XL U2301 ( .A0(n273), .A1(n1776), .B0(n2314), .B1(n209), .Y(n529) );
  OAI22XL U2302 ( .A0(n273), .A1(n1778), .B0(n2314), .B1(n1777), .Y(n528) );
  OAI22XL U2303 ( .A0(n273), .A1(n1779), .B0(n2314), .B1(n203), .Y(n527) );
  OAI22XL U2304 ( .A0(n273), .A1(n964), .B0(n2314), .B1(n107), .Y(n526) );
  OAI22XL U2305 ( .A0(n273), .A1(n1780), .B0(n2314), .B1(n227), .Y(n525) );
  OAI22XL U2306 ( .A0(n273), .A1(n175), .B0(n2314), .B1(n211), .Y(n524) );
  OAI22XL U2307 ( .A0(n273), .A1(n787), .B0(n2314), .B1(n230), .Y(n523) );
  OAI22XL U2308 ( .A0(n273), .A1(n174), .B0(n2314), .B1(n229), .Y(n522) );
  OA22X1 U2309 ( .A0(n1782), .A1(n1965), .B0(n212), .B1(n1785), .Y(n1787) );
  AO21X1 U2310 ( .A0(n1803), .A1(n1801), .B0(n1798), .Y(n1804) );
  OAI21XL U2311 ( .A0(n1801), .A1(n1798), .B0(n1800), .Y(n1799) );
  OAI21XL U2312 ( .A0(n1813), .A1(n1812), .B0(n1816), .Y(n1814) );
  OA21XL U2313 ( .A0(n1960), .A1(n1826), .B0(n110), .Y(n1833) );
  OAI2BB1X1 U2314 ( .A0N(n1837), .A1N(n1830), .B0(n1952), .Y(n1832) );
  OAI21XL U2315 ( .A0(n1830), .A1(n1829), .B0(n1833), .Y(n1831) );
  OR2X1 U2316 ( .A(n120), .B(n1835), .Y(n1843) );
  OAI2BB1X1 U2317 ( .A0N(n1843), .A1N(n1841), .B0(n1955), .Y(n1844) );
  OAI21XL U2318 ( .A0(n1841), .A1(n1838), .B0(n1840), .Y(n1839) );
  OR2X1 U2319 ( .A(n1847), .B(n1846), .Y(n1855) );
  OAI2BB1X1 U2320 ( .A0N(n1855), .A1N(n1852), .B0(n1946), .Y(n1848) );
  OAI2BB1X1 U2321 ( .A0N(n1857), .A1N(n1860), .B0(n1954), .Y(n1862) );
  OAI21XL U2322 ( .A0(n1860), .A1(n1859), .B0(n1863), .Y(n1861) );
  OR2X1 U2323 ( .A(n1869), .B(n1864), .Y(n1873) );
  OAI2BB1X1 U2324 ( .A0N(n1873), .A1N(n1868), .B0(n1949), .Y(n1870) );
  OA21XL U2325 ( .A0(n1949), .A1(n1872), .B0(n1870), .Y(n1881) );
  OAI2BB1X1 U2326 ( .A0N(n1875), .A1N(n1878), .B0(n1956), .Y(n1880) );
  OAI21XL U2327 ( .A0(n1878), .A1(n1877), .B0(n1881), .Y(n1879) );
  OR2X1 U2328 ( .A(n118), .B(n1882), .Y(n1888) );
  OAI2BB1X1 U2329 ( .A0N(n1888), .A1N(n1886), .B0(n1948), .Y(n1889) );
  OA21XL U2330 ( .A0(n1948), .A1(n1890), .B0(n1889), .Y(n1897) );
  OAI2BB1X1 U2331 ( .A0N(n1900), .A1N(n1894), .B0(n1947), .Y(n1896) );
  OAI21XL U2332 ( .A0(n1894), .A1(n1893), .B0(n1897), .Y(n1895) );
  OR2X1 U2333 ( .A(n121), .B(n1898), .Y(n1905) );
  OAI2BB1X1 U2334 ( .A0N(n1905), .A1N(n1903), .B0(n1908), .Y(n1906) );
  OAI21XL U2335 ( .A0(n1903), .A1(n1953), .B0(n1902), .Y(n1901) );
  OR2X1 U2336 ( .A(n1910), .B(n1909), .Y(n1921) );
  OAI2BB1X1 U2337 ( .A0N(n1921), .A1N(n1915), .B0(n1911), .Y(n1917) );
  OAI21XL U2338 ( .A0(n1915), .A1(n1914), .B0(n1918), .Y(n1916) );
  OR2X1 U2339 ( .A(n1919), .B(n1926), .Y(n1927) );
  OAI2BB1X1 U2340 ( .A0N(n1927), .A1N(n1925), .B0(n2120), .Y(n1928) );
  OAI21XL U2341 ( .A0(n1922), .A1(n1925), .B0(n1924), .Y(n1923) );
  OA21XL U2342 ( .A0(n1935), .A1(n1934), .B0(n1936), .Y(n1943) );
  OAI31XL U2343 ( .A0(n1940), .A1(n1939), .A2(n1938), .B0(n1937), .Y(n1941) );
  AOI2BB1X1 U2344 ( .A0N(n1945), .A1N(n234), .B0(n1941), .Y(n1942) );
  OAI22XL U2345 ( .A0(n1945), .A1(n1944), .B0(n1943), .B1(n1942), .Y(n2118) );
  OAI21XL U2346 ( .A0(curr_photo_size[1]), .A1(n1968), .B0(curr_photo_size[0]), 
        .Y(n2116) );
  AOI2BB1X1 U2347 ( .A0N(n1972), .A1N(n212), .B0(n2114), .Y(n1978) );
  OA21XL U2348 ( .A0(n1974), .A1(n213), .B0(n1976), .Y(n1977) );
  AOI222XL U2349 ( .A0(n1999), .A1(n1991), .B0(n1999), .B1(n182), .C0(n1991), 
        .C1(n1990), .Y(n1986) );
  AOI2BB2X1 U2350 ( .B0(n1987), .B1(n1993), .A0N(n1987), .A1N(n1986), .Y(n1998) );
  OAI21XL U2351 ( .A0(n1995), .A1(n1994), .B0(n1993), .Y(n1996) );
  OAI21XL U2352 ( .A0(work_cntr[15]), .A1(n2012), .B0(n1998), .Y(n2000) );
  OAI21XL U2353 ( .A0(work_cntr[14]), .A1(n2014), .B0(n2011), .Y(n2002) );
  NOR3BXL U2354 ( .AN(n2012), .B(n2011), .C(n2009), .Y(n2005) );
  NAND3BX1 U2355 ( .AN(n2005), .B(n2006), .C(n2014), .Y(n2022) );
  OAI21XL U2356 ( .A0(n2009), .A1(n2011), .B0(n2012), .Y(n2010) );
  OAI21XL U2357 ( .A0(work_cntr[13]), .A1(n2027), .B0(n2013), .Y(n2016) );
  OAI21XL U2358 ( .A0(work_cntr[12]), .A1(n2030), .B0(n2021), .Y(n2018) );
  OAI21XL U2359 ( .A0(work_cntr[11]), .A1(n2044), .B0(n2029), .Y(n2032) );
  OAI21XL U2360 ( .A0(work_cntr[10]), .A1(n2047), .B0(n2037), .Y(n2034) );
  OAI21XL U2361 ( .A0(work_cntr[9]), .A1(n2063), .B0(n2046), .Y(n2049) );
  OAI21XL U2362 ( .A0(work_cntr[8]), .A1(n2066), .B0(n2054), .Y(n2051) );
  OAI21XL U2363 ( .A0(work_cntr[7]), .A1(n2079), .B0(n2065), .Y(n2068) );
  OAI21XL U2364 ( .A0(work_cntr[6]), .A1(n2082), .B0(n2073), .Y(n2070) );
  OAI21XL U2365 ( .A0(work_cntr[5]), .A1(n2092), .B0(n2081), .Y(n2084) );
  OAI21XL U2366 ( .A0(work_cntr[4]), .A1(n2102), .B0(n2089), .Y(n2086) );
  AOI2BB2X1 U2367 ( .B0(n2088), .B1(n2087), .A0N(n2088), .A1N(n2086), .Y(n2095) );
  AOI2BB1X1 U2368 ( .A0N(n2095), .A1N(n2102), .B0(n2098), .Y(n2106) );
  AOI2BB2X1 U2369 ( .B0(N2062), .B1(n2107), .A0N(N2062), .A1N(n2107), .Y(n2109) );
  AO21X1 U2370 ( .A0(n2111), .A1(N2061), .B0(N85), .Y(n2108) );
  OAI21XL U2371 ( .A0(n2111), .A1(N2061), .B0(n2110), .Y(n2113) );
  OAI22XL U2372 ( .A0(n2114), .A1(n2113), .B0(n2112), .B1(n2323), .Y(n2115) );
  OAI22XL U2373 ( .A0(n2277), .A1(sftr_n[1]), .B0(n2116), .B1(n2115), .Y(n2117) );
  AO21X1 U2374 ( .A0(n2118), .A1(n716), .B0(n2117), .Y(n2287) );
  OR2X1 U2375 ( .A(next_work_cntr[17]), .B(n2131), .Y(n2130) );
  OAI21XL U2376 ( .A0(n2120), .A1(n179), .B0(next_work_cntr[1]), .Y(n2121) );
  AOI2BB2X1 U2377 ( .B0(next_work_cntr[19]), .B1(n2129), .A0N(
        next_work_cntr[19]), .A1N(n2129), .Y(n2136) );
  AOI2BB2X1 U2378 ( .B0(next_work_cntr[16]), .B1(n2132), .A0N(n2132), .A1N(
        next_work_cntr[16]), .Y(n2134) );
  AOI2BB2X1 U2379 ( .B0(n2140), .B1(next_work_cntr[15]), .A0N(n2140), .A1N(
        next_work_cntr[15]), .Y(n2143) );
  AOI2BB1X1 U2380 ( .A0N(n2153), .A1N(n2150), .B0(n2149), .Y(n2152) );
  AOI2BB1X1 U2381 ( .A0N(n2161), .A1N(n2157), .B0(n2156), .Y(n2160) );
  NAND3BX1 U2382 ( .AN(n2175), .B(n2166), .C(n2169), .Y(n2171) );
  AOI2BB2X1 U2383 ( .B0(n2169), .B1(n2168), .A0N(n2169), .A1N(n2168), .Y(n2172) );
  AOI2BB2X1 U2384 ( .B0(n2186), .B1(n2185), .A0N(n2186), .A1N(n2185), .Y(n2189) );
  AOI2BB2X1 U2385 ( .B0(n2192), .B1(n2191), .A0N(n2192), .A1N(n2191), .Y(n2202) );
  AOI2BB2X1 U2386 ( .B0(n2197), .B1(n2196), .A0N(n2197), .A1N(n2196), .Y(n2198) );
  OAI31XL U2387 ( .A0(n2202), .A1(n2204), .A2(n2219), .B0(n2198), .Y(n2200) );
  AOI2BB1X1 U2388 ( .A0N(n2206), .A1N(n2200), .B0(n2199), .Y(n2201) );
  OAI21XL U2389 ( .A0(n2219), .A1(n2208), .B0(n2207), .Y(n2213) );
  AOI2BB2X1 U2390 ( .B0(next_work_cntr[6]), .B1(n2217), .A0N(n2217), .A1N(
        next_work_cntr[6]), .Y(n2223) );
  OAI21XL U2391 ( .A0(n2220), .A1(n2229), .B0(n2219), .Y(n2218) );
  OAI21XL U2392 ( .A0(n2229), .A1(n2228), .B0(n2231), .Y(n2230) );
  AOI2BB2X1 U2393 ( .B0(n2241), .B1(n2240), .A0N(n2241), .A1N(n2240), .Y(n2242) );
  OAI21XL U2394 ( .A0(n2246), .A1(n2244), .B0(n2245), .Y(n2243) );
  OA21XL U2395 ( .A0(n2260), .A1(n2259), .B0(n2258), .Y(n2275) );
  AOI2BB2X1 U2396 ( .B0(n2262), .B1(n2261), .A0N(n2262), .A1N(n2261), .Y(n2273) );
  OAI2BB1X1 U2397 ( .A0N(n2265), .A1N(n2264), .B0(n2263), .Y(n2266) );
  OAI22XL U2398 ( .A0(n2277), .A1(n2276), .B0(n2275), .B1(n2274), .Y(n2286) );
  OAI31XL U2399 ( .A0(n2316), .A1(si_sel), .A2(n2315), .B0(n2283), .Y(n2285)
         );
  OAI2BB1X1 U2400 ( .A0N(n2287), .A1N(n690), .B0(n2291), .Y(next_en_si) );
  OAI2BB2XL U2401 ( .B0(cr_read_cntr[4]), .B1(n2296), .A0N(cr_read_cntr[4]), 
        .A1N(n2295), .Y(n495) );
  OA21XL U2402 ( .A0(cr_read_cntr[6]), .A1(n2300), .B0(n2301), .Y(n493) );
  OAI22XL U2403 ( .A0(n240), .A1(photo_num[1]), .B0(n188), .B1(photo_num[0]), 
        .Y(n2317) );
  AOI2BB2X1 U2404 ( .B0(n2333), .B1(n2332), .A0N(n2331), .A1N(sftr_n[1]), .Y(
        n2335) );
endmodule


module DPA ( clk, reset, IM_A, IM_Q, IM_D, IM_WEN, CR_A, CR_Q );
  output [19:0] IM_A;
  input [23:0] IM_Q;
  output [23:0] IM_D;
  output [8:0] CR_A;
  input [12:0] CR_Q;
  input clk, reset;
  output IM_WEN;
  wire   n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, im_d_w_19,
         im_d_w_18, im_d_w_9, im_d_w_8, en_si, en_init_time, en_fb_addr,
         en_photo_num, en_curr_photo_size, en_so, si_sel, init_time_mux_sel,
         \sftr_n[1] , \data_path/si_w[0] , \data_path/si_w[1] ,
         \data_path/si_w[2] , \data_path/si_w[3] , \data_path/si_w[4] ,
         \data_path/si_w[5] , \data_path/si_w[6] , \data_path/si_w[7] ,
         \data_path/si_w[8] , \data_path/si_w[9] , \data_path/si_w[10] ,
         \data_path/si_w[11] , \data_path/si_w[12] , \data_path/si_w[13] ,
         \data_path/si_w[14] , \data_path/si_w[15] , \data_path/si_w[16] ,
         \data_path/si_w[17] , \data_path/si_w[18] , \data_path/si_w[19] ,
         \data_path/si_w[20] , \data_path/si_w[21] , \data_path/si_w[22] ,
         \data_path/si_w[23] , n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n141, n144, n145, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, \intadd_0/CI , \intadd_0/SUM[6] ,
         \intadd_0/SUM[5] , \intadd_0/SUM[4] , \intadd_0/SUM[3] ,
         \intadd_0/SUM[2] , \intadd_0/SUM[1] , \intadd_0/SUM[0] ,
         \intadd_0/n7 , \intadd_0/n6 , \intadd_0/n5 , \intadd_0/n4 ,
         \intadd_0/n3 , \intadd_0/n2 , \intadd_0/n1 , \intadd_1/CI ,
         \intadd_1/SUM[6] , \intadd_1/SUM[5] , \intadd_1/SUM[4] ,
         \intadd_1/SUM[3] , \intadd_1/SUM[2] , \intadd_1/SUM[1] ,
         \intadd_1/SUM[0] , \intadd_1/n7 , \intadd_1/n6 , \intadd_1/n5 ,
         \intadd_1/n4 , \intadd_1/n3 , \intadd_1/n2 , \intadd_1/n1 ,
         \intadd_2/CI , \intadd_2/SUM[6] , \intadd_2/SUM[5] ,
         \intadd_2/SUM[4] , \intadd_2/SUM[3] , \intadd_2/SUM[2] ,
         \intadd_2/SUM[1] , \intadd_2/SUM[0] , \intadd_2/n7 , \intadd_2/n6 ,
         \intadd_2/n5 , \intadd_2/n4 , \intadd_2/n3 , \intadd_2/n2 ,
         \intadd_2/n1 , n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n442, n444, n446, n448, n450, n452, n454, n456, n458, n460, n462,
         n463, n464, n465, n466, n467, n468, n469, n471, n473, n475, n477,
         n480, n482, n484, n486, n488, n490, n492, n494, n496, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n757;
  wire   [29:28] im_d_w;
  wire   [23:0] curr_time;
  wire   [19:0] fb_addr;
  wire   [1:0] photo_num;
  wire   [19:0] curr_photo_addr;
  wire   [1:0] curr_photo_size;
  wire   [1:0] so_mux_sel;
  wire   [3:0] expand_sel;
  wire   SYNOPSYS_UNCONNECTED__0;

  CONT ctrl_logic ( .clk(clk), .reset(reset), .im_wen_n(IM_WEN), .cr_a(CR_A), 
        .curr_time(curr_time), .fb_addr(fb_addr), .photo_num(photo_num), 
        .curr_photo_addr(curr_photo_addr), .curr_photo_size(curr_photo_size), 
        .en_si(en_si), .en_init_time(en_init_time), .en_fb_addr(en_fb_addr), 
        .en_photo_num(en_photo_num), .en_curr_photo_addr(n467), 
        .en_curr_photo_size(en_curr_photo_size), .en_so(en_so), .si_sel(si_sel), .init_time_mux_sel(init_time_mux_sel), .sftr_n({\sftr_n[1] , 
        SYNOPSYS_UNCONNECTED__0}), .so_mux_sel(so_mux_sel), .expand_sel({
        expand_sel[3], n464, expand_sel[1:0]}), .\im_a[19]_BAR (n758), 
        .\im_a[18]_BAR (n759), .\im_a[17]_BAR (n760), .\im_a[16]_BAR (n761), 
        .\im_a[15]_BAR (n762), .\im_a[14]_BAR (n763), .\im_a[13]_BAR (n764), 
        .\im_a[12]_BAR (n765), .\im_a[11]_BAR (n766), .\im_a[10]_BAR (n767), 
        .\im_a[9]_BAR (n768), .\im_a[8]_BAR (n769), .\im_a[7]_BAR (n770), 
        .\im_a[6]_BAR (n771), .\im_a[5]_BAR (n772), .\im_a[4]_BAR (n773), 
        .\im_a[3]_BAR (n774), .\im_a[2]_BAR (n775), .\im_a[1]_BAR (n776), 
        .\im_a[0]_BAR (n777) );
  ADDFXL \intadd_0/U3  ( .A(n779), .B(\data_path/si_w[22] ), .CI(\intadd_0/n3 ), .CO(\intadd_0/n2 ), .S(\intadd_0/SUM[5] ) );
  ADDFXL \intadd_1/U3  ( .A(IM_D[14]), .B(\data_path/si_w[14] ), .CI(
        \intadd_1/n3 ), .CO(\intadd_1/n2 ), .S(\intadd_1/SUM[5] ) );
  ADDFXL \intadd_2/U3  ( .A(IM_D[6]), .B(\data_path/si_w[6] ), .CI(
        \intadd_2/n3 ), .CO(\intadd_2/n2 ), .S(\intadd_2/SUM[5] ) );
  DFFSX1 \data_path/si_reg/q_reg[2]  ( .D(n314), .CK(clk), .SN(n22), .Q(n509), 
        .QN(\data_path/si_w[2] ) );
  DFFSX1 \data_path/si_reg/q_reg[4]  ( .D(n313), .CK(clk), .SN(n463), .Q(n508), 
        .QN(\data_path/si_w[4] ) );
  DFFSX1 \data_path/si_reg/q_reg[1]  ( .D(n315), .CK(clk), .SN(n463), .Q(n503), 
        .QN(\data_path/si_w[1] ) );
  DFFSX1 \data_path/si_reg/q_reg[8]  ( .D(n312), .CK(clk), .SN(n462), .Q(n499), 
        .QN(\data_path/si_w[8] ) );
  DFFSX1 \data_path/init_time_reg/q_reg[1]  ( .D(n145), .CK(clk), .SN(n463), 
        .Q(n652), .QN(curr_time[1]) );
  ADDFXL \intadd_1/U2  ( .A(IM_D[15]), .B(\data_path/si_w[15] ), .CI(
        \intadd_1/n2 ), .CO(\intadd_1/n1 ), .S(\intadd_1/SUM[6] ) );
  ADDFXL \intadd_0/U2  ( .A(n778), .B(\data_path/si_w[23] ), .CI(\intadd_0/n2 ), .CO(\intadd_0/n1 ), .S(\intadd_0/SUM[6] ) );
  ADDFXL \intadd_2/U2  ( .A(IM_D[7]), .B(\data_path/si_w[7] ), .CI(
        \intadd_2/n2 ), .CO(\intadd_2/n1 ), .S(\intadd_2/SUM[6] ) );
  ADDFXL \intadd_1/U8  ( .A(n787), .B(\data_path/si_w[9] ), .CI(\intadd_1/CI ), 
        .CO(\intadd_1/n7 ), .S(\intadd_1/SUM[0] ) );
  ADDFXL \intadd_1/U7  ( .A(n786), .B(\data_path/si_w[10] ), .CI(\intadd_1/n7 ), .CO(\intadd_1/n6 ), .S(\intadd_1/SUM[1] ) );
  ADDFXL \intadd_1/U6  ( .A(n785), .B(\data_path/si_w[11] ), .CI(\intadd_1/n6 ), .CO(\intadd_1/n5 ), .S(\intadd_1/SUM[2] ) );
  ADDFXL \intadd_1/U5  ( .A(IM_D[12]), .B(\data_path/si_w[12] ), .CI(
        \intadd_1/n5 ), .CO(\intadd_1/n4 ), .S(\intadd_1/SUM[3] ) );
  ADDFXL \intadd_1/U4  ( .A(IM_D[13]), .B(\data_path/si_w[13] ), .CI(
        \intadd_1/n4 ), .CO(\intadd_1/n3 ), .S(\intadd_1/SUM[4] ) );
  ADDFXL \intadd_0/U8  ( .A(IM_D[17]), .B(\data_path/si_w[17] ), .CI(
        \intadd_0/CI ), .CO(\intadd_0/n7 ), .S(\intadd_0/SUM[0] ) );
  ADDFXL \intadd_0/U7  ( .A(IM_D[18]), .B(\data_path/si_w[18] ), .CI(
        \intadd_0/n7 ), .CO(\intadd_0/n6 ), .S(\intadd_0/SUM[1] ) );
  ADDFXL \intadd_0/U6  ( .A(n782), .B(\data_path/si_w[19] ), .CI(\intadd_0/n6 ), .CO(\intadd_0/n5 ), .S(\intadd_0/SUM[2] ) );
  ADDFXL \intadd_0/U5  ( .A(n781), .B(\data_path/si_w[20] ), .CI(\intadd_0/n5 ), .CO(\intadd_0/n4 ), .S(\intadd_0/SUM[3] ) );
  ADDFXL \intadd_0/U4  ( .A(n780), .B(\data_path/si_w[21] ), .CI(\intadd_0/n4 ), .CO(\intadd_0/n3 ), .S(\intadd_0/SUM[4] ) );
  ADDFXL \intadd_2/U8  ( .A(IM_D[1]), .B(\data_path/si_w[1] ), .CI(
        \intadd_2/CI ), .CO(\intadd_2/n7 ), .S(\intadd_2/SUM[0] ) );
  ADDFXL \intadd_2/U7  ( .A(IM_D[2]), .B(\data_path/si_w[2] ), .CI(
        \intadd_2/n7 ), .CO(\intadd_2/n6 ), .S(\intadd_2/SUM[1] ) );
  ADDFXL \intadd_2/U6  ( .A(IM_D[3]), .B(\data_path/si_w[3] ), .CI(
        \intadd_2/n6 ), .CO(\intadd_2/n5 ), .S(\intadd_2/SUM[2] ) );
  ADDFXL \intadd_2/U5  ( .A(IM_D[4]), .B(\data_path/si_w[4] ), .CI(
        \intadd_2/n5 ), .CO(\intadd_2/n4 ), .S(\intadd_2/SUM[3] ) );
  ADDFXL \intadd_2/U4  ( .A(IM_D[5]), .B(\data_path/si_w[5] ), .CI(
        \intadd_2/n4 ), .CO(\intadd_2/n3 ), .S(\intadd_2/SUM[4] ) );
  DFFRX2 \data_path/si_reg/q_reg[0]  ( .D(n417), .CK(clk), .RN(n462), .Q(
        \data_path/si_w[0] ), .QN(n514) );
  DFFSX2 \data_path/init_time_reg/q_reg[4]  ( .D(n141), .CK(clk), .SN(n462), 
        .QN(curr_time[4]) );
  DFFRX2 \data_path/init_time_reg/q_reg[17]  ( .D(n322), .CK(clk), .RN(n22), 
        .Q(curr_time[17]), .QN(n505) );
  DFFRX2 \data_path/init_time_reg/q_reg[12]  ( .D(n327), .CK(clk), .RN(n463), 
        .Q(curr_time[12]), .QN(n518) );
  DFFSX2 \data_path/init_time_reg/q_reg[2]  ( .D(n144), .CK(clk), .SN(n463), 
        .QN(curr_time[2]) );
  DFFRX2 \data_path/init_time_reg/q_reg[19]  ( .D(n320), .CK(clk), .RN(n462), 
        .Q(curr_time[19]), .QN(n531) );
  DFFRX2 \data_path/init_time_reg/q_reg[15]  ( .D(n324), .CK(clk), .RN(n462), 
        .Q(curr_time[15]) );
  DFFRX2 \data_path/init_time_reg/q_reg[9]  ( .D(n330), .CK(clk), .RN(n463), 
        .Q(curr_time[9]), .QN(n529) );
  DFFRX2 \data_path/init_time_reg/q_reg[11]  ( .D(n328), .CK(clk), .RN(n462), 
        .Q(curr_time[11]), .QN(n500) );
  DFFRX2 \data_path/init_time_reg/q_reg[7]  ( .D(n332), .CK(clk), .RN(n462), 
        .Q(curr_time[7]) );
  DFFRX2 \data_path/init_time_reg/q_reg[6]  ( .D(n333), .CK(clk), .RN(n22), 
        .Q(curr_time[6]) );
  DFFRX2 \data_path/init_time_reg/q_reg[14]  ( .D(n325), .CK(clk), .RN(n22), 
        .Q(curr_time[14]) );
  DFFRX1 \data_path/photo_num_reg/q_reg[0]  ( .D(n367), .CK(clk), .RN(n462), 
        .Q(photo_num[0]) );
  DFFRX1 \data_path/si_reg/q_reg[16]  ( .D(n418), .CK(clk), .RN(n22), .Q(
        \data_path/si_w[16] ) );
  DFFRX1 \data_path/si_reg/q_reg[11]  ( .D(n396), .CK(clk), .RN(n463), .Q(
        \data_path/si_w[11] ), .QN(n714) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[16]  ( .D(n12), .CK(clk), .RN(n462), .Q(
        fb_addr[16]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[0]  ( .D(n415), .CK(clk), .RN(
        n22), .Q(curr_photo_addr[0]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[2]  ( .D(n17), .CK(clk), .RN(
        n463), .Q(curr_photo_addr[2]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[15]  ( .D(n382), .CK(clk), .RN(
        n462), .Q(curr_photo_addr[15]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[14]  ( .D(n385), .CK(clk), .RN(
        n22), .Q(curr_photo_addr[14]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[4]  ( .D(n15), .CK(clk), .RN(
        n463), .Q(curr_photo_addr[4]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[19]  ( .D(n373), .CK(clk), .RN(
        n462), .Q(curr_photo_addr[19]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[18]  ( .D(n376), .CK(clk), .RN(
        n22), .Q(curr_photo_addr[18]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[17]  ( .D(n379), .CK(clk), .RN(
        n463), .Q(curr_photo_addr[17]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[9]  ( .D(n400), .CK(clk), .RN(
        n462), .Q(curr_photo_addr[9]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[6]  ( .D(n406), .CK(clk), .RN(
        n22), .Q(curr_photo_addr[6]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[12]  ( .D(n391), .CK(clk), .RN(
        n463), .Q(curr_photo_addr[12]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[10]  ( .D(n397), .CK(clk), .RN(
        n462), .Q(curr_photo_addr[10]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[5]  ( .D(n409), .CK(clk), .RN(
        n22), .Q(curr_photo_addr[5]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[1]  ( .D(n19), .CK(clk), .RN(
        n463), .Q(curr_photo_addr[1]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[8]  ( .D(n13), .CK(clk), .RN(
        n462), .Q(curr_photo_addr[8]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[7]  ( .D(n403), .CK(clk), .RN(
        n22), .Q(curr_photo_addr[7]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[3]  ( .D(n412), .CK(clk), .RN(
        n463), .Q(curr_photo_addr[3]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[13]  ( .D(n388), .CK(clk), .RN(
        n462), .Q(curr_photo_addr[13]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[11]  ( .D(n394), .CK(clk), .RN(
        n22), .Q(curr_photo_addr[11]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[16]  ( .D(n11), .CK(clk), .RN(
        n463), .Q(curr_photo_addr[16]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[6]  ( .D(n407), .CK(clk), .RN(n462), .Q(
        fb_addr[6]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[5]  ( .D(n410), .CK(clk), .RN(n22), .Q(
        fb_addr[5]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[0]  ( .D(n416), .CK(clk), .RN(n463), .Q(
        fb_addr[0]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[9]  ( .D(n401), .CK(clk), .RN(n462), .Q(
        fb_addr[9]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[7]  ( .D(n404), .CK(clk), .RN(n22), .Q(
        fb_addr[7]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[13]  ( .D(n389), .CK(clk), .RN(n463), 
        .Q(fb_addr[13]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[19]  ( .D(n374), .CK(clk), .RN(n462), 
        .Q(fb_addr[19]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[18]  ( .D(n377), .CK(clk), .RN(n22), .Q(
        fb_addr[18]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[17]  ( .D(n380), .CK(clk), .RN(n463), 
        .Q(fb_addr[17]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[15]  ( .D(n383), .CK(clk), .RN(n462), 
        .Q(fb_addr[15]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[14]  ( .D(n386), .CK(clk), .RN(n22), .Q(
        fb_addr[14]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[12]  ( .D(n392), .CK(clk), .RN(n463), 
        .Q(fb_addr[12]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[11]  ( .D(n395), .CK(clk), .RN(n462), 
        .Q(fb_addr[11]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[10]  ( .D(n398), .CK(clk), .RN(n22), .Q(
        fb_addr[10]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[4]  ( .D(n16), .CK(clk), .RN(n463), .Q(
        fb_addr[4]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[2]  ( .D(n18), .CK(clk), .RN(n462), .Q(
        fb_addr[2]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[1]  ( .D(n20), .CK(clk), .RN(n22), .Q(
        fb_addr[1]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[8]  ( .D(n14), .CK(clk), .RN(n463), .Q(
        fb_addr[8]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[3]  ( .D(n413), .CK(clk), .RN(n462), .Q(
        fb_addr[3]) );
  DFFRX1 \data_path/init_time_reg/q_reg[5]  ( .D(n334), .CK(clk), .RN(n22), 
        .Q(curr_time[5]) );
  DFFRX1 \data_path/init_time_reg/q_reg[8]  ( .D(n331), .CK(clk), .RN(n463), 
        .Q(curr_time[8]) );
  DFFRX1 \data_path/so_reg/q_reg[29]  ( .D(n337), .CK(clk), .RN(n462), .Q(
        im_d_w[29]) );
  DFFRX1 \data_path/so_reg/q_reg[19]  ( .D(n347), .CK(clk), .RN(n22), .Q(
        im_d_w_19) );
  DFFRX1 \data_path/so_reg/q_reg[9]  ( .D(n357), .CK(clk), .RN(n463), .Q(
        im_d_w_9) );
  DFFRX1 \data_path/so_reg/q_reg[17]  ( .D(n349), .CK(clk), .RN(n462), .QN(
        n494) );
  DFFRX1 \data_path/so_reg/q_reg[7]  ( .D(n359), .CK(clk), .RN(n22), .QN(n496)
         );
  DFFRX1 \data_path/so_reg/q_reg[1]  ( .D(n365), .CK(clk), .RN(n463), .QN(n477) );
  DFFRX1 \data_path/so_reg/q_reg[22]  ( .D(n344), .CK(clk), .RN(n462), .Q(n783) );
  DFFRX1 \data_path/so_reg/q_reg[21]  ( .D(n345), .CK(clk), .RN(n22), .QN(n475) );
  DFFRX1 \data_path/so_reg/q_reg[16]  ( .D(n350), .CK(clk), .RN(n463), .QN(
        n473) );
  DFFRX1 \data_path/so_reg/q_reg[15]  ( .D(n351), .CK(clk), .RN(n462), .QN(
        n484) );
  DFFRX1 \data_path/so_reg/q_reg[14]  ( .D(n352), .CK(clk), .RN(n22), .QN(n486) );
  DFFRX1 \data_path/so_reg/q_reg[6]  ( .D(n360), .CK(clk), .RN(n463), .QN(n492) );
  DFFRX1 \data_path/so_reg/q_reg[5]  ( .D(n361), .CK(clk), .RN(n462), .QN(n490) );
  DFFRX1 \data_path/so_reg/q_reg[4]  ( .D(n362), .CK(clk), .RN(n22), .QN(n488)
         );
  DFFRX1 \data_path/so_reg/q_reg[3]  ( .D(n363), .CK(clk), .RN(n463), .QN(n482) );
  DFFRX1 \data_path/so_reg/q_reg[2]  ( .D(n364), .CK(clk), .RN(n462), .QN(n480) );
  DFFRX1 \data_path/si_reg/q_reg[23]  ( .D(n369), .CK(clk), .RN(n22), .Q(
        \data_path/si_w[23] ), .QN(n512) );
  DFFRX1 \data_path/si_reg/q_reg[22]  ( .D(n370), .CK(clk), .RN(n463), .Q(
        \data_path/si_w[22] ), .QN(n511) );
  DFFRX1 \data_path/si_reg/q_reg[21]  ( .D(n371), .CK(clk), .RN(n462), .Q(
        \data_path/si_w[21] ), .QN(n510) );
  DFFRX1 \data_path/si_reg/q_reg[20]  ( .D(n372), .CK(clk), .RN(n22), .Q(
        \data_path/si_w[20] ), .QN(n532) );
  DFFRX1 \data_path/si_reg/q_reg[19]  ( .D(n375), .CK(clk), .RN(n463), .Q(
        \data_path/si_w[19] ), .QN(n526) );
  DFFRX1 \data_path/si_reg/q_reg[18]  ( .D(n378), .CK(clk), .RN(n462), .Q(
        \data_path/si_w[18] ), .QN(n524) );
  DFFRX1 \data_path/si_reg/q_reg[17]  ( .D(n381), .CK(clk), .RN(n22), .Q(
        \data_path/si_w[17] ), .QN(n525) );
  DFFRX1 \data_path/si_reg/q_reg[15]  ( .D(n384), .CK(clk), .RN(n463), .Q(
        \data_path/si_w[15] ), .QN(n523) );
  DFFRX1 \data_path/si_reg/q_reg[14]  ( .D(n387), .CK(clk), .RN(n462), .Q(
        \data_path/si_w[14] ), .QN(n527) );
  DFFRX1 \data_path/si_reg/q_reg[13]  ( .D(n390), .CK(clk), .RN(n22), .Q(
        \data_path/si_w[13] ), .QN(n506) );
  DFFRX1 \data_path/photo_num_reg/q_reg[1]  ( .D(n21), .CK(clk), .RN(n463), 
        .Q(photo_num[1]), .QN(n10) );
  DFFRX1 \data_path/si_reg/q_reg[12]  ( .D(n393), .CK(clk), .RN(n462), .Q(
        \data_path/si_w[12] ), .QN(n520) );
  DFFRX1 \data_path/si_reg/q_reg[10]  ( .D(n399), .CK(clk), .RN(n22), .Q(
        \data_path/si_w[10] ), .QN(n498) );
  DFFRX1 \data_path/si_reg/q_reg[9]  ( .D(n402), .CK(clk), .RN(n463), .Q(
        \data_path/si_w[9] ), .QN(n521) );
  DFFRX1 \data_path/si_reg/q_reg[7]  ( .D(n405), .CK(clk), .RN(n462), .Q(
        \data_path/si_w[7] ), .QN(n517) );
  DFFRX1 \data_path/si_reg/q_reg[6]  ( .D(n408), .CK(clk), .RN(n22), .Q(
        \data_path/si_w[6] ), .QN(n522) );
  DFFRX1 \data_path/si_reg/q_reg[5]  ( .D(n411), .CK(clk), .RN(n463), .Q(
        \data_path/si_w[5] ), .QN(n507) );
  DFFRX1 \data_path/si_reg/q_reg[3]  ( .D(n414), .CK(clk), .RN(n462), .Q(
        \data_path/si_w[3] ), .QN(n516) );
  DFFRX1 \data_path/curr_photo_size_reg/q_reg[1]  ( .D(n23), .CK(clk), .RN(n22), .Q(curr_photo_size[1]), .QN(n535) );
  DFFRX1 \data_path/curr_photo_size_reg/q_reg[0]  ( .D(n368), .CK(clk), .RN(
        n463), .Q(curr_photo_size[0]), .QN(n513) );
  DFFRX1 \data_path/init_time_reg/q_reg[16]  ( .D(n323), .CK(clk), .RN(n462), 
        .Q(curr_time[16]), .QN(n501) );
  DFFRX1 \data_path/init_time_reg/q_reg[0]  ( .D(n336), .CK(clk), .RN(n22), 
        .Q(curr_time[0]), .QN(n515) );
  DFFRX1 \data_path/init_time_reg/q_reg[18]  ( .D(n321), .CK(clk), .RN(n463), 
        .Q(curr_time[18]), .QN(n519) );
  DFFRX1 \data_path/init_time_reg/q_reg[23]  ( .D(n316), .CK(clk), .RN(n462), 
        .Q(curr_time[23]), .QN(n502) );
  DFFRX1 \data_path/init_time_reg/q_reg[22]  ( .D(n317), .CK(clk), .RN(n22), 
        .Q(curr_time[22]), .QN(n530) );
  DFFRX1 \data_path/init_time_reg/q_reg[21]  ( .D(n318), .CK(clk), .RN(n463), 
        .Q(curr_time[21]), .QN(n534) );
  DFFRX1 \data_path/init_time_reg/q_reg[13]  ( .D(n326), .CK(clk), .RN(n462), 
        .Q(curr_time[13]), .QN(n533) );
  DFFRX1 \data_path/init_time_reg/q_reg[3]  ( .D(n335), .CK(clk), .RN(n22), 
        .Q(curr_time[3]), .QN(n528) );
  DFFRX1 \data_path/init_time_reg/q_reg[10]  ( .D(n329), .CK(clk), .RN(n463), 
        .Q(curr_time[10]), .QN(n504) );
  DFFRX1 \data_path/so_reg/q_reg[28]  ( .D(n338), .CK(clk), .RN(n462), .Q(
        im_d_w[28]), .QN(n537) );
  DFFRX1 \data_path/so_reg/q_reg[18]  ( .D(n348), .CK(clk), .RN(n22), .Q(
        im_d_w_18), .QN(n538) );
  DFFRX1 \data_path/so_reg/q_reg[8]  ( .D(n358), .CK(clk), .RN(n463), .Q(
        im_d_w_8), .QN(n536) );
  DFFRX1 \data_path/so_reg/q_reg[27]  ( .D(n339), .CK(clk), .RN(n462), .Q(n778), .QN(n454) );
  DFFRX1 \data_path/so_reg/q_reg[20]  ( .D(n346), .CK(clk), .RN(n22), .Q(n784), 
        .QN(n460) );
  DFFRX1 \data_path/so_reg/q_reg[10]  ( .D(n356), .CK(clk), .RN(n463), .Q(n788), .QN(n458) );
  DFFRX1 \data_path/so_reg/q_reg[0]  ( .D(n366), .CK(clk), .RN(n462), .Q(n789), 
        .QN(n456) );
  DFFRX1 \data_path/so_reg/q_reg[26]  ( .D(n340), .CK(clk), .RN(n22), .Q(n779), 
        .QN(n452) );
  DFFRX1 \data_path/so_reg/q_reg[25]  ( .D(n341), .CK(clk), .RN(n463), .Q(n780), .QN(n450) );
  DFFRX1 \data_path/so_reg/q_reg[24]  ( .D(n342), .CK(clk), .RN(n462), .Q(n781), .QN(n448) );
  DFFRX1 \data_path/so_reg/q_reg[23]  ( .D(n343), .CK(clk), .RN(n22), .Q(n782), 
        .QN(n446) );
  DFFRX1 \data_path/so_reg/q_reg[13]  ( .D(n353), .CK(clk), .RN(n463), .Q(n785), .QN(n444) );
  DFFRX1 \data_path/so_reg/q_reg[12]  ( .D(n354), .CK(clk), .RN(n22), .Q(n786), 
        .QN(n442) );
  DFFRX1 \data_path/so_reg/q_reg[11]  ( .D(n355), .CK(clk), .RN(n463), .Q(n787), .QN(n440) );
  DFFRX2 \data_path/init_time_reg/q_reg[20]  ( .D(n319), .CK(clk), .RN(n22), 
        .Q(curr_time[20]) );
  BUFX4 U435 ( .A(n733), .Y(n542) );
  CLKBUFX3 U436 ( .A(n734), .Y(n543) );
  AO22X1 U437 ( .A0(n539), .A1(\intadd_0/SUM[2] ), .B0(\intadd_0/SUM[1] ), 
        .B1(n540), .Y(n421) );
  AOI211XL U438 ( .A0(IM_D[17]), .A1(n730), .B0(n637), .C0(n421), .Y(n422) );
  NAND2X1 U439 ( .A(\intadd_0/SUM[0] ), .B(n541), .Y(n423) );
  OAI211XL U440 ( .A0(n465), .A1(n525), .B0(n422), .C0(n423), .Y(n345) );
  AO22X1 U441 ( .A0(n539), .A1(\intadd_0/SUM[3] ), .B0(\intadd_0/SUM[2] ), 
        .B1(n540), .Y(n424) );
  AOI211XL U442 ( .A0(IM_D[18]), .A1(n730), .B0(n637), .C0(n424), .Y(n425) );
  NAND2XL U443 ( .A(\intadd_0/SUM[1] ), .B(n541), .Y(n426) );
  OAI211XL U444 ( .A0(n465), .A1(n524), .B0(n425), .C0(n426), .Y(n344) );
  AO22X1 U445 ( .A0(n539), .A1(\intadd_2/SUM[2] ), .B0(n540), .B1(
        \intadd_2/SUM[1] ), .Y(n427) );
  AOI211X1 U446 ( .A0(IM_D[1]), .A1(n730), .B0(n637), .C0(n427), .Y(n428) );
  NAND2X1 U447 ( .A(\intadd_2/SUM[0] ), .B(n541), .Y(n429) );
  OAI211XL U448 ( .A0(n465), .A1(n503), .B0(n428), .C0(n429), .Y(n365) );
  NOR4X1 U449 ( .A(n468), .B(\data_path/si_w[17] ), .C(\data_path/si_w[18] ), 
        .D(\data_path/si_w[19] ), .Y(n430) );
  NOR4X1 U450 ( .A(\data_path/si_w[1] ), .B(\data_path/si_w[2] ), .C(
        \data_path/si_w[15] ), .D(\data_path/si_w[23] ), .Y(n431) );
  NOR4X1 U451 ( .A(\data_path/si_w[20] ), .B(\data_path/si_w[14] ), .C(
        \data_path/si_w[21] ), .D(\data_path/si_w[22] ), .Y(n432) );
  AND4X1 U452 ( .A(n431), .B(n432), .C(n520), .D(en_curr_photo_size), .Y(n433)
         );
  AND4X1 U453 ( .A(n499), .B(n430), .C(n506), .D(n433), .Y(n551) );
  NOR2X1 U454 ( .A(n642), .B(n703), .Y(n434) );
  OAI2BB2XL U455 ( .B0(n517), .B1(n465), .A0N(\intadd_2/SUM[6] ), .A1N(n541), 
        .Y(n435) );
  AOI211X1 U456 ( .A0(IM_D[7]), .A1(n730), .B0(n434), .C0(n435), .Y(n436) );
  OAI211X1 U457 ( .A0(n729), .A1(n597), .B0(n647), .C0(n436), .Y(n359) );
  NOR2X1 U458 ( .A(n642), .B(n732), .Y(n437) );
  OAI2BB2XL U459 ( .B0(n465), .B1(n523), .A0N(\intadd_1/SUM[6] ), .A1N(n541), 
        .Y(n438) );
  AOI211X1 U460 ( .A0(IM_D[15]), .A1(n730), .B0(n437), .C0(n438), .Y(n439) );
  OAI211X1 U461 ( .A0(n729), .A1(n728), .B0(n647), .C0(n439), .Y(n349) );
  INVX16 U462 ( .A(n440), .Y(IM_D[9]) );
  INVX16 U463 ( .A(n442), .Y(IM_D[10]) );
  INVX16 U464 ( .A(n444), .Y(IM_D[11]) );
  INVX16 U465 ( .A(n446), .Y(IM_D[19]) );
  INVX16 U466 ( .A(n448), .Y(IM_D[20]) );
  INVX16 U467 ( .A(n450), .Y(IM_D[21]) );
  INVX16 U468 ( .A(n452), .Y(IM_D[22]) );
  INVX16 U469 ( .A(n454), .Y(IM_D[23]) );
  INVX16 U470 ( .A(n456), .Y(IM_D[0]) );
  INVX16 U471 ( .A(n458), .Y(IM_D[8]) );
  INVX16 U472 ( .A(n460), .Y(IM_D[16]) );
  INVX8 U473 ( .A(reset), .Y(n462) );
  INVX8 U474 ( .A(reset), .Y(n463) );
  INVX8 U475 ( .A(reset), .Y(n22) );
  NOR2X2 U476 ( .A(expand_sel[1]), .B(expand_sel[0]), .Y(n572) );
  CLKBUFX4 U477 ( .A(n644), .Y(n465) );
  NOR2X1 U478 ( .A(n660), .B(n662), .Y(n668) );
  INVX1 U479 ( .A(en_fb_addr), .Y(n547) );
  INVX6 U480 ( .A(n544), .Y(n466) );
  INVX4 U481 ( .A(en_so), .Y(n730) );
  INVX2 U482 ( .A(en_si), .Y(n734) );
  NAND3BXL U483 ( .AN(so_mux_sel[0]), .B(en_so), .C(n556), .Y(n644) );
  AOI211X1 U484 ( .A0(n690), .A1(curr_time[20]), .B0(n679), .C0(n678), .Y(n681) );
  INVX1 U485 ( .A(n467), .Y(n544) );
  NOR2X1 U486 ( .A(si_sel), .B(n543), .Y(n733) );
  INVX16 U487 ( .A(n484), .Y(IM_D[13]) );
  BUFX16 U488 ( .A(n783), .Y(IM_D[18]) );
  CLKBUFX2 U489 ( .A(\data_path/si_w[16] ), .Y(n468) );
  NAND2X1 U490 ( .A(n712), .B(n711), .Y(n722) );
  NOR2X1 U491 ( .A(n504), .B(n710), .Y(n711) );
  NOR2X1 U492 ( .A(n528), .B(n660), .Y(n663) );
  NAND2X1 U493 ( .A(curr_time[2]), .B(n657), .Y(n660) );
  NOR2X1 U494 ( .A(n701), .B(n726), .Y(n705) );
  NOR2X1 U495 ( .A(curr_time[8]), .B(n717), .Y(n701) );
  CLKINVX1 U496 ( .A(n651), .Y(n662) );
  NOR2X1 U497 ( .A(n673), .B(n666), .Y(n651) );
  NOR2X1 U498 ( .A(n501), .B(n688), .Y(n683) );
  NAND2X1 U499 ( .A(en_init_time), .B(n681), .Y(n688) );
  AOI211X1 U500 ( .A0(curr_time[13]), .A1(n672), .B0(curr_time[15]), .C0(
        curr_time[14]), .Y(n679) );
  AOI211X1 U501 ( .A0(n649), .A1(curr_time[5]), .B0(curr_time[6]), .C0(
        curr_time[7]), .Y(n671) );
  OAI21X1 U502 ( .A0(curr_time[16]), .A1(n689), .B0(n724), .Y(n684) );
  CLKINVX1 U503 ( .A(n681), .Y(n689) );
  AOI211X1 U504 ( .A0(curr_time[2]), .A1(n657), .B0(n673), .C0(n666), .Y(n658)
         );
  OAI21X1 U505 ( .A0(n690), .A1(n689), .B0(n724), .Y(n693) );
  NOR2BX1 U506 ( .AN(n690), .B(n688), .Y(n692) );
  NOR3X2 U507 ( .A(n505), .B(n501), .C(n519), .Y(n690) );
  OAI21X1 U508 ( .A0(\intadd_0/n1 ), .A1(im_d_w[28]), .B0(n641), .Y(n695) );
  NAND2X1 U509 ( .A(\intadd_0/n1 ), .B(im_d_w[28]), .Y(n641) );
  OAI31X1 U510 ( .A0(n563), .A1(n562), .A2(n561), .B0(expand_sel[3]), .Y(n577)
         );
  CLKINVX1 U511 ( .A(n539), .Y(n642) );
  BUFX4 U512 ( .A(n632), .Y(n539) );
  BUFX4 U513 ( .A(n638), .Y(n540) );
  INVX3 U514 ( .A(n547), .Y(n546) );
  CLKINVX1 U515 ( .A(n738), .Y(n469) );
  INVX16 U516 ( .A(n469), .Y(IM_A[0]) );
  INVX16 U517 ( .A(n776), .Y(IM_A[1]) );
  INVX16 U518 ( .A(n775), .Y(IM_A[2]) );
  INVX16 U519 ( .A(n774), .Y(IM_A[3]) );
  INVX16 U520 ( .A(n773), .Y(IM_A[4]) );
  INVX16 U521 ( .A(n772), .Y(IM_A[5]) );
  INVX16 U522 ( .A(n771), .Y(IM_A[6]) );
  INVX16 U523 ( .A(n770), .Y(IM_A[7]) );
  INVX16 U524 ( .A(n769), .Y(IM_A[8]) );
  INVX16 U525 ( .A(n768), .Y(IM_A[9]) );
  INVX16 U526 ( .A(n767), .Y(IM_A[10]) );
  INVX16 U527 ( .A(n766), .Y(IM_A[11]) );
  INVX16 U528 ( .A(n765), .Y(IM_A[12]) );
  INVX16 U529 ( .A(n764), .Y(IM_A[13]) );
  INVX16 U530 ( .A(n763), .Y(IM_A[14]) );
  INVX16 U531 ( .A(n762), .Y(IM_A[15]) );
  INVX16 U532 ( .A(n761), .Y(IM_A[16]) );
  INVX16 U533 ( .A(n760), .Y(IM_A[17]) );
  INVX16 U534 ( .A(n759), .Y(IM_A[18]) );
  CLKINVX1 U535 ( .A(n757), .Y(n471) );
  INVX16 U536 ( .A(n471), .Y(IM_A[19]) );
  INVX16 U537 ( .A(n473), .Y(IM_D[14]) );
  INVX16 U538 ( .A(n475), .Y(IM_D[17]) );
  INVX16 U539 ( .A(n477), .Y(IM_D[1]) );
  INVX16 U540 ( .A(n480), .Y(IM_D[2]) );
  INVX16 U541 ( .A(n482), .Y(IM_D[3]) );
  INVX16 U542 ( .A(n486), .Y(IM_D[12]) );
  INVX16 U543 ( .A(n488), .Y(IM_D[4]) );
  INVX16 U544 ( .A(n490), .Y(IM_D[5]) );
  INVX16 U545 ( .A(n492), .Y(IM_D[6]) );
  INVX16 U546 ( .A(n494), .Y(IM_D[15]) );
  INVX16 U547 ( .A(n496), .Y(IM_D[7]) );
  NAND2X1 U548 ( .A(n556), .B(so_mux_sel[0]), .Y(n621) );
  OAI21X1 U549 ( .A0(\intadd_2/n1 ), .A1(im_d_w_8), .B0(n596), .Y(n597) );
  NAND2X1 U550 ( .A(\intadd_2/n1 ), .B(im_d_w_8), .Y(n596) );
  OAI21X1 U551 ( .A0(\intadd_1/n1 ), .A1(im_d_w_18), .B0(n620), .Y(n728) );
  NAND2X1 U552 ( .A(\intadd_1/n1 ), .B(im_d_w_18), .Y(n620) );
  NAND2X1 U553 ( .A(expand_sel[0]), .B(n569), .Y(n570) );
  CLKINVX1 U554 ( .A(expand_sel[1]), .Y(n569) );
  NOR2X1 U555 ( .A(\data_path/si_w[4] ), .B(n549), .Y(n552) );
  NAND4X1 U556 ( .A(n498), .B(n714), .C(n507), .D(n522), .Y(n549) );
  NOR2BX1 U557 ( .AN(init_time_mux_sel), .B(n671), .Y(n677) );
  NAND2X1 U558 ( .A(n671), .B(init_time_mux_sel), .Y(n666) );
  CLKINVX1 U559 ( .A(n712), .Y(n717) );
  NOR2X1 U560 ( .A(n675), .B(n673), .Y(n712) );
  NAND2XL U561 ( .A(IM_D[14]), .B(n730), .Y(n618) );
  NOR2X1 U562 ( .A(curr_time[2]), .B(n657), .Y(n655) );
  NOR2X2 U563 ( .A(n652), .B(n515), .Y(n657) );
  BUFX4 U564 ( .A(n643), .Y(n541) );
  NOR2XL U565 ( .A(n730), .B(n621), .Y(n643) );
  INVX3 U566 ( .A(n727), .Y(n725) );
  NOR2X4 U567 ( .A(init_time_mux_sel), .B(n673), .Y(n727) );
  INVX4 U568 ( .A(n647), .Y(n637) );
  NAND4X2 U569 ( .A(so_mux_sel[1]), .B(n578), .C(n577), .D(n576), .Y(n647) );
  NOR2BX2 U570 ( .AN(n675), .B(n726), .Y(n724) );
  NAND2X2 U571 ( .A(en_init_time), .B(n666), .Y(n726) );
  NAND2XL U572 ( .A(n779), .B(n730), .Y(n639) );
  AOI211XL U573 ( .A0(n778), .A1(n730), .B0(n646), .C0(n645), .Y(n648) );
  INVX3 U574 ( .A(n547), .Y(n545) );
  AOI22XL U575 ( .A0(\data_path/si_w[8] ), .A1(n599), .B0(n788), .B1(n598), 
        .Y(n600) );
  AOI22XL U576 ( .A0(\data_path/si_w[0] ), .A1(n558), .B0(n789), .B1(n557), 
        .Y(n579) );
  AOI22XL U577 ( .A0(n468), .A1(n623), .B0(n784), .B1(n622), .Y(n624) );
  INVXL U578 ( .A(en_photo_num), .Y(n736) );
  OAI211XL U579 ( .A0(en_curr_photo_size), .A1(n513), .B0(n554), .C0(n737), 
        .Y(n368) );
  NAND4XL U580 ( .A(\data_path/si_w[7] ), .B(n552), .C(n551), .D(n550), .Y(
        n554) );
  NOR3XL U581 ( .A(\data_path/si_w[9] ), .B(\data_path/si_w[0] ), .C(
        \data_path/si_w[3] ), .Y(n550) );
  INVXL U582 ( .A(n698), .Y(n411) );
  INVXL U583 ( .A(n704), .Y(n402) );
  INVXL U584 ( .A(n699), .Y(n408) );
  INVXL U585 ( .A(n548), .Y(n417) );
  INVXL U586 ( .A(n697), .Y(n414) );
  INVXL U587 ( .A(n709), .Y(n399) );
  INVXL U588 ( .A(n715), .Y(n396) );
  INVXL U589 ( .A(n721), .Y(n393) );
  INVXL U590 ( .A(n700), .Y(n405) );
  NAND4XL U591 ( .A(n553), .B(n552), .C(n551), .D(n517), .Y(n737) );
  INVXL U592 ( .A(n655), .Y(n656) );
  AOI211XL U593 ( .A0(curr_time[4]), .A1(n673), .B0(n665), .C0(n664), .Y(n141)
         );
  NOR2XL U594 ( .A(n725), .B(n508), .Y(n664) );
  AOI211XL U595 ( .A0(curr_time[4]), .A1(n663), .B0(n662), .C0(n661), .Y(n665)
         );
  NOR2XL U596 ( .A(curr_time[4]), .B(n663), .Y(n661) );
  NOR2XL U597 ( .A(n654), .B(n653), .Y(n145) );
  AOI211XL U598 ( .A0(n652), .A1(n515), .B0(n657), .C0(n662), .Y(n654) );
  INVXL U599 ( .A(n670), .Y(n334) );
  INVXL U600 ( .A(n667), .Y(n669) );
  OAI32XL U601 ( .A0(n528), .A1(n658), .A2(n673), .B0(n668), .B1(curr_time[3]), 
        .Y(n659) );
  NAND2XL U602 ( .A(curr_time[12]), .B(curr_time[11]), .Y(n723) );
  AOI21XL U603 ( .A0(curr_time[8]), .A1(n726), .B0(n701), .Y(n674) );
  AOI22XL U604 ( .A0(curr_time[12]), .A1(n718), .B0(n727), .B1(
        \data_path/si_w[12] ), .Y(n719) );
  AOI22XL U605 ( .A0(curr_time[10]), .A1(n706), .B0(\data_path/si_w[10] ), 
        .B1(n727), .Y(n707) );
  NAND2XL U606 ( .A(curr_time[8]), .B(n712), .Y(n708) );
  OAI211XL U607 ( .A0(n725), .A1(n524), .B0(n687), .C0(n686), .Y(n321) );
  NOR2XL U608 ( .A(n689), .B(curr_time[17]), .Y(n685) );
  NAND3XL U609 ( .A(curr_time[17]), .B(n683), .C(n519), .Y(n687) );
  INVXL U610 ( .A(n694), .Y(n319) );
  CLKINVX2 U611 ( .A(en_init_time), .Y(n673) );
  NAND2XL U612 ( .A(n677), .B(n679), .Y(n675) );
  NAND3XL U613 ( .A(n677), .B(n676), .C(n502), .Y(n678) );
  AOI211XL U614 ( .A0(curr_time[20]), .A1(curr_time[19]), .B0(curr_time[21]), 
        .C0(curr_time[22]), .Y(n676) );
  NOR2XL U615 ( .A(n655), .B(n667), .Y(n649) );
  NAND2XL U616 ( .A(curr_time[4]), .B(curr_time[3]), .Y(n667) );
  AOI211XL U617 ( .A0(n504), .A1(n710), .B0(n518), .C0(n500), .Y(n672) );
  NAND2XL U618 ( .A(curr_time[9]), .B(curr_time[8]), .Y(n710) );
  OAI211XL U619 ( .A0(n729), .A1(n695), .B0(n648), .C0(n647), .Y(n339) );
  NOR2XL U620 ( .A(n642), .B(n696), .Y(n646) );
  NAND3XL U621 ( .A(n625), .B(n624), .C(n647), .Y(n346) );
  OAI21XL U622 ( .A0(n784), .A1(n731), .B0(n465), .Y(n623) );
  AOI22XL U623 ( .A0(n539), .A1(\intadd_0/SUM[1] ), .B0(n540), .B1(
        \intadd_0/SUM[0] ), .Y(n625) );
  NAND3XL U624 ( .A(n601), .B(n600), .C(n647), .Y(n356) );
  OAI21XL U625 ( .A0(n788), .A1(n731), .B0(n465), .Y(n599) );
  AOI22XL U626 ( .A0(n539), .A1(\intadd_1/SUM[1] ), .B0(n540), .B1(
        \intadd_1/SUM[0] ), .Y(n601) );
  NAND3XL U627 ( .A(n580), .B(n579), .C(n647), .Y(n366) );
  OAI21XL U628 ( .A0(n789), .A1(n731), .B0(n465), .Y(n558) );
  INVX3 U629 ( .A(n541), .Y(n731) );
  AOI22XL U630 ( .A0(n539), .A1(\intadd_2/SUM[1] ), .B0(n540), .B1(
        \intadd_2/SUM[0] ), .Y(n580) );
  OAI211XL U631 ( .A0(n465), .A1(n521), .B0(n604), .C0(n603), .Y(n355) );
  NAND2XL U632 ( .A(n541), .B(\intadd_1/SUM[0] ), .Y(n603) );
  AOI211XL U633 ( .A0(n540), .A1(\intadd_1/SUM[1] ), .B0(n637), .C0(n602), .Y(
        n604) );
  OAI211XL U634 ( .A0(n465), .A1(n507), .B0(n592), .C0(n591), .Y(n361) );
  NAND2XL U635 ( .A(n541), .B(\intadd_2/SUM[4] ), .Y(n591) );
  AOI211XL U636 ( .A0(n540), .A1(\intadd_2/SUM[5] ), .B0(n637), .C0(n590), .Y(
        n592) );
  OAI211XL U637 ( .A0(n465), .A1(n714), .B0(n610), .C0(n609), .Y(n353) );
  NAND2XL U638 ( .A(n541), .B(\intadd_1/SUM[2] ), .Y(n609) );
  AOI211XL U639 ( .A0(n540), .A1(\intadd_1/SUM[3] ), .B0(n637), .C0(n608), .Y(
        n610) );
  OAI211XL U640 ( .A0(n465), .A1(n498), .B0(n607), .C0(n606), .Y(n354) );
  NAND2XL U641 ( .A(n541), .B(\intadd_1/SUM[1] ), .Y(n606) );
  AOI211XL U642 ( .A0(n540), .A1(\intadd_1/SUM[2] ), .B0(n637), .C0(n605), .Y(
        n607) );
  OAI211XL U643 ( .A0(n506), .A1(n465), .B0(n616), .C0(n615), .Y(n351) );
  NAND2XL U644 ( .A(n541), .B(\intadd_1/SUM[4] ), .Y(n615) );
  AOI211XL U645 ( .A0(n540), .A1(\intadd_1/SUM[5] ), .B0(n637), .C0(n614), .Y(
        n616) );
  OAI211XL U646 ( .A0(n465), .A1(n516), .B0(n586), .C0(n585), .Y(n363) );
  NAND2XL U647 ( .A(n541), .B(\intadd_2/SUM[2] ), .Y(n585) );
  AOI211XL U648 ( .A0(n540), .A1(\intadd_2/SUM[3] ), .B0(n637), .C0(n584), .Y(
        n586) );
  OAI211XL U649 ( .A0(n465), .A1(n508), .B0(n589), .C0(n588), .Y(n362) );
  NAND2XL U650 ( .A(n541), .B(\intadd_2/SUM[3] ), .Y(n588) );
  AOI211XL U651 ( .A0(n540), .A1(\intadd_2/SUM[4] ), .B0(n637), .C0(n587), .Y(
        n589) );
  OAI211XL U652 ( .A0(n465), .A1(n532), .B0(n631), .C0(n630), .Y(n342) );
  NAND2XL U653 ( .A(n541), .B(\intadd_0/SUM[3] ), .Y(n630) );
  AOI211XL U654 ( .A0(n540), .A1(\intadd_0/SUM[4] ), .B0(n637), .C0(n629), .Y(
        n631) );
  OAI211XL U655 ( .A0(n465), .A1(n520), .B0(n613), .C0(n612), .Y(n352) );
  NAND2XL U656 ( .A(n541), .B(\intadd_1/SUM[3] ), .Y(n612) );
  AOI211XL U657 ( .A0(n540), .A1(\intadd_1/SUM[4] ), .B0(n637), .C0(n611), .Y(
        n613) );
  OAI211XL U658 ( .A0(n465), .A1(n526), .B0(n628), .C0(n627), .Y(n343) );
  NAND2XL U659 ( .A(n541), .B(\intadd_0/SUM[2] ), .Y(n627) );
  AOI211XL U660 ( .A0(n540), .A1(\intadd_0/SUM[3] ), .B0(n637), .C0(n626), .Y(
        n628) );
  OAI211XL U661 ( .A0(n510), .A1(n465), .B0(n635), .C0(n634), .Y(n341) );
  NAND2XL U662 ( .A(n541), .B(\intadd_0/SUM[4] ), .Y(n634) );
  AOI211XL U663 ( .A0(n540), .A1(\intadd_0/SUM[5] ), .B0(n637), .C0(n633), .Y(
        n635) );
  OAI211XL U664 ( .A0(n465), .A1(n509), .B0(n583), .C0(n582), .Y(n364) );
  NAND2XL U665 ( .A(n541), .B(\intadd_2/SUM[1] ), .Y(n582) );
  AOI211XL U666 ( .A0(n540), .A1(\intadd_2/SUM[2] ), .B0(n637), .C0(n581), .Y(
        n583) );
  OAI211XL U667 ( .A0(n597), .A1(n642), .B0(n595), .C0(n594), .Y(n360) );
  NAND2X1 U668 ( .A(IM_D[6]), .B(n730), .Y(n594) );
  AOI211XL U669 ( .A0(n540), .A1(\intadd_2/SUM[6] ), .B0(n637), .C0(n593), .Y(
        n595) );
  NOR2BXL U670 ( .AN(n789), .B(n514), .Y(\intadd_2/CI ) );
  OAI211XL U671 ( .A0(n695), .A1(n642), .B0(n640), .C0(n639), .Y(n340) );
  AOI211XL U672 ( .A0(n540), .A1(\intadd_0/SUM[6] ), .B0(n637), .C0(n636), .Y(
        n640) );
  AND2XL U673 ( .A(n468), .B(n784), .Y(\intadd_0/CI ) );
  OAI211XL U674 ( .A0(n728), .A1(n642), .B0(n619), .C0(n618), .Y(n350) );
  AOI211XL U675 ( .A0(n540), .A1(\intadd_1/SUM[6] ), .B0(n637), .C0(n617), .Y(
        n619) );
  INVXL U676 ( .A(so_mux_sel[1]), .Y(n556) );
  INVXL U677 ( .A(expand_sel[3]), .Y(n573) );
  AOI211XL U678 ( .A0(n572), .A1(\data_path/si_w[12] ), .B0(n464), .C0(n571), 
        .Y(n574) );
  AOI211XL U679 ( .A0(n572), .A1(\data_path/si_w[8] ), .B0(n566), .C0(n565), 
        .Y(n575) );
  AOI211XL U680 ( .A0(n572), .A1(\data_path/si_w[4] ), .B0(n464), .C0(n560), 
        .Y(n561) );
  INVXL U681 ( .A(expand_sel[0]), .Y(n567) );
  NOR2XL U682 ( .A(\data_path/si_w[0] ), .B(n566), .Y(n562) );
  NOR2XL U683 ( .A(n572), .B(n566), .Y(n563) );
  INVXL U684 ( .A(n464), .Y(n566) );
  NOR2XL U685 ( .A(so_mux_sel[0]), .B(n730), .Y(n578) );
  NOR2BXL U686 ( .AN(\sftr_n[1] ), .B(n555), .Y(n632) );
  NAND3XL U687 ( .A(so_mux_sel[1]), .B(so_mux_sel[0]), .C(en_so), .Y(n555) );
  NOR2BXL U688 ( .AN(n788), .B(n499), .Y(\intadd_1/CI ) );
  INVXL U689 ( .A(n777), .Y(n738) );
  INVXL U690 ( .A(n758), .Y(n757) );
  AOI222XL U691 ( .A0(n543), .A1(\data_path/si_w[8] ), .B0(n542), .B1(IM_Q[8]), 
        .C0(n720), .C1(CR_Q[8]), .Y(n312) );
  AOI222XL U692 ( .A0(n543), .A1(\data_path/si_w[4] ), .B0(n542), .B1(IM_Q[4]), 
        .C0(n720), .C1(CR_Q[4]), .Y(n313) );
  AOI222XL U693 ( .A0(n734), .A1(\data_path/si_w[2] ), .B0(n542), .B1(IM_Q[2]), 
        .C0(n720), .C1(CR_Q[2]), .Y(n314) );
  AOI222XL U694 ( .A0(n543), .A1(\data_path/si_w[1] ), .B0(n720), .B1(CR_Q[1]), 
        .C0(IM_Q[1]), .C1(n542), .Y(n315) );
  OAI22XL U695 ( .A0(en_photo_num), .A1(n10), .B0(n736), .B1(n735), .Y(n21) );
  AOI222XL U696 ( .A0(n543), .A1(\data_path/si_w[5] ), .B0(n542), .B1(IM_Q[5]), 
        .C0(n720), .C1(CR_Q[5]), .Y(n698) );
  AOI222XL U697 ( .A0(n543), .A1(\data_path/si_w[9] ), .B0(n542), .B1(IM_Q[9]), 
        .C0(n720), .C1(CR_Q[9]), .Y(n704) );
  AOI222XL U698 ( .A0(n543), .A1(\data_path/si_w[6] ), .B0(n542), .B1(IM_Q[6]), 
        .C0(n720), .C1(CR_Q[6]), .Y(n699) );
  AOI222XL U699 ( .A0(n543), .A1(\data_path/si_w[0] ), .B0(n542), .B1(IM_Q[0]), 
        .C0(n720), .C1(CR_Q[0]), .Y(n548) );
  AOI222XL U700 ( .A0(n543), .A1(\data_path/si_w[3] ), .B0(n542), .B1(IM_Q[3]), 
        .C0(n720), .C1(CR_Q[3]), .Y(n697) );
  AOI222XL U701 ( .A0(n543), .A1(\data_path/si_w[10] ), .B0(n542), .B1(
        IM_Q[10]), .C0(n720), .C1(CR_Q[10]), .Y(n709) );
  AOI222XL U702 ( .A0(n543), .A1(\data_path/si_w[11] ), .B0(n542), .B1(
        IM_Q[11]), .C0(n720), .C1(CR_Q[11]), .Y(n715) );
  AOI222XL U703 ( .A0(n543), .A1(\data_path/si_w[12] ), .B0(n542), .B1(
        IM_Q[12]), .C0(n720), .C1(CR_Q[12]), .Y(n721) );
  AOI222XL U704 ( .A0(n543), .A1(\data_path/si_w[7] ), .B0(n542), .B1(IM_Q[7]), 
        .C0(n720), .C1(CR_Q[7]), .Y(n700) );
  AND2X2 U705 ( .A(si_sel), .B(en_si), .Y(n720) );
  NOR3XL U706 ( .A(\data_path/si_w[0] ), .B(\data_path/si_w[3] ), .C(n521), 
        .Y(n553) );
  AOI222XL U707 ( .A0(n673), .A1(curr_time[2]), .B0(n727), .B1(
        \data_path/si_w[2] ), .C0(n656), .C1(n658), .Y(n144) );
  AOI222XL U708 ( .A0(\data_path/si_w[5] ), .A1(n727), .B0(curr_time[5]), .B1(
        n726), .C0(n669), .C1(n668), .Y(n670) );
  OAI222XL U709 ( .A0(n506), .A1(n725), .B0(n533), .B1(n724), .C0(n723), .C1(
        n722), .Y(n326) );
  OAI21XL U710 ( .A0(n716), .A1(n500), .B0(n713), .Y(n328) );
  OAI31XL U711 ( .A0(curr_time[12]), .A1(n500), .A2(n722), .B0(n719), .Y(n327)
         );
  OAI31XL U712 ( .A0(curr_time[10]), .A1(n529), .A2(n708), .B0(n707), .Y(n329)
         );
  AOI222XL U713 ( .A0(n693), .A1(curr_time[20]), .B0(curr_time[19]), .B1(n692), 
        .C0(n727), .C1(\data_path/si_w[20] ), .Y(n694) );
  CLKINVX1 U714 ( .A(n540), .Y(n729) );
  NOR2X1 U715 ( .A(\sftr_n[1] ), .B(n555), .Y(n638) );
  AO22X1 U716 ( .A0(n468), .A1(n734), .B0(n542), .B1(IM_Q[16]), .Y(n418) );
  AOI2BB2X1 U717 ( .B0(n546), .B1(n514), .A0N(en_fb_addr), .A1N(fb_addr[0]), 
        .Y(n416) );
  AOI2BB2X1 U718 ( .B0(n466), .B1(n514), .A0N(n466), .A1N(curr_photo_addr[0]), 
        .Y(n415) );
  AOI2BB2X1 U719 ( .B0(n546), .B1(n516), .A0N(n545), .A1N(fb_addr[3]), .Y(n413) );
  AOI2BB2X1 U720 ( .B0(n466), .B1(n516), .A0N(n466), .A1N(curr_photo_addr[3]), 
        .Y(n412) );
  AOI2BB2X1 U721 ( .B0(n546), .B1(n507), .A0N(en_fb_addr), .A1N(fb_addr[5]), 
        .Y(n410) );
  AOI2BB2X1 U722 ( .B0(n466), .B1(n507), .A0N(n466), .A1N(curr_photo_addr[5]), 
        .Y(n409) );
  AOI2BB2X1 U723 ( .B0(n546), .B1(n522), .A0N(en_fb_addr), .A1N(fb_addr[6]), 
        .Y(n407) );
  AOI2BB2X1 U724 ( .B0(n466), .B1(n522), .A0N(n466), .A1N(curr_photo_addr[6]), 
        .Y(n406) );
  AOI2BB2X1 U725 ( .B0(n546), .B1(n517), .A0N(n546), .A1N(fb_addr[7]), .Y(n404) );
  AOI2BB2X1 U726 ( .B0(n466), .B1(n517), .A0N(n466), .A1N(curr_photo_addr[7]), 
        .Y(n403) );
  AOI2BB2X1 U727 ( .B0(en_photo_num), .B1(\data_path/si_w[0] ), .A0N(
        en_photo_num), .A1N(photo_num[0]), .Y(n367) );
  OAI21XL U728 ( .A0(\data_path/si_w[0] ), .A1(n621), .B0(en_so), .Y(n557) );
  OAI22XL U729 ( .A0(expand_sel[0]), .A1(\data_path/si_w[2] ), .B0(n567), .B1(
        \data_path/si_w[1] ), .Y(n559) );
  OAI22XL U730 ( .A0(n569), .A1(n559), .B0(n516), .B1(n570), .Y(n560) );
  OAI22XL U731 ( .A0(expand_sel[0]), .A1(\data_path/si_w[6] ), .B0(n567), .B1(
        \data_path/si_w[5] ), .Y(n564) );
  OAI22XL U732 ( .A0(n569), .A1(n564), .B0(n570), .B1(n517), .Y(n565) );
  OAI22XL U733 ( .A0(expand_sel[0]), .A1(\data_path/si_w[10] ), .B0(n567), 
        .B1(\data_path/si_w[9] ), .Y(n568) );
  OAI22XL U734 ( .A0(n714), .A1(n570), .B0(n569), .B1(n568), .Y(n571) );
  OAI21XL U735 ( .A0(n575), .A1(n574), .B0(n573), .Y(n576) );
  AO22X1 U736 ( .A0(\intadd_2/SUM[3] ), .A1(n539), .B0(IM_D[2]), .B1(n730), 
        .Y(n581) );
  AO22X1 U737 ( .A0(\intadd_2/SUM[4] ), .A1(n539), .B0(IM_D[3]), .B1(n730), 
        .Y(n584) );
  AO22X1 U738 ( .A0(\intadd_2/SUM[5] ), .A1(n539), .B0(IM_D[4]), .B1(n730), 
        .Y(n587) );
  AO22X1 U739 ( .A0(\intadd_2/SUM[6] ), .A1(n539), .B0(IM_D[5]), .B1(n730), 
        .Y(n590) );
  OAI2BB2XL U740 ( .B0(n522), .B1(n465), .A0N(n541), .A1N(\intadd_2/SUM[5] ), 
        .Y(n593) );
  AOI2BB2X1 U741 ( .B0(im_d_w_9), .B1(n596), .A0N(im_d_w_9), .A1N(n596), .Y(
        n703) );
  OAI222XL U742 ( .A0(n703), .A1(n729), .B0(n536), .B1(en_so), .C0(n597), .C1(
        n731), .Y(n358) );
  OAI21XL U743 ( .A0(\data_path/si_w[8] ), .A1(n621), .B0(en_so), .Y(n598) );
  AO22X1 U744 ( .A0(\intadd_1/SUM[2] ), .A1(n539), .B0(n787), .B1(n730), .Y(
        n602) );
  AO22X1 U745 ( .A0(\intadd_1/SUM[3] ), .A1(n539), .B0(n786), .B1(n730), .Y(
        n605) );
  AO22X1 U746 ( .A0(\intadd_1/SUM[4] ), .A1(n539), .B0(n785), .B1(n730), .Y(
        n608) );
  AO22X1 U747 ( .A0(\intadd_1/SUM[5] ), .A1(n539), .B0(IM_D[12]), .B1(n730), 
        .Y(n611) );
  AO22X1 U748 ( .A0(\intadd_1/SUM[6] ), .A1(n539), .B0(IM_D[13]), .B1(n730), 
        .Y(n614) );
  OAI2BB2XL U749 ( .B0(n465), .B1(n527), .A0N(n541), .A1N(\intadd_1/SUM[5] ), 
        .Y(n617) );
  AOI2BB2X1 U750 ( .B0(im_d_w_19), .B1(n620), .A0N(im_d_w_19), .A1N(n620), .Y(
        n732) );
  OAI21XL U751 ( .A0(n468), .A1(n621), .B0(en_so), .Y(n622) );
  AO22X1 U752 ( .A0(\intadd_0/SUM[4] ), .A1(n539), .B0(n782), .B1(n730), .Y(
        n626) );
  AO22X1 U753 ( .A0(\intadd_0/SUM[5] ), .A1(n539), .B0(n781), .B1(n730), .Y(
        n629) );
  AO22X1 U754 ( .A0(\intadd_0/SUM[6] ), .A1(n539), .B0(n780), .B1(n730), .Y(
        n633) );
  OAI2BB2XL U755 ( .B0(n465), .B1(n511), .A0N(n541), .A1N(\intadd_0/SUM[5] ), 
        .Y(n636) );
  AOI2BB2X1 U756 ( .B0(im_d_w[29]), .B1(n641), .A0N(im_d_w[29]), .A1N(n641), 
        .Y(n696) );
  OAI2BB2XL U757 ( .B0(n465), .B1(n512), .A0N(n541), .A1N(\intadd_0/SUM[6] ), 
        .Y(n645) );
  OAI22XL U758 ( .A0(curr_time[0]), .A1(n651), .B0(n515), .B1(n673), .Y(n650)
         );
  OAI21XL U759 ( .A0(n725), .A1(n514), .B0(n650), .Y(n336) );
  OAI22XL U760 ( .A0(en_init_time), .A1(n652), .B0(n725), .B1(n503), .Y(n653)
         );
  OAI21XL U761 ( .A0(n725), .A1(n516), .B0(n659), .Y(n335) );
  AO22X1 U762 ( .A0(n727), .A1(\data_path/si_w[6] ), .B0(n673), .B1(
        curr_time[6]), .Y(n333) );
  AO22X1 U763 ( .A0(n727), .A1(\data_path/si_w[7] ), .B0(n673), .B1(
        curr_time[7]), .Y(n332) );
  OAI21XL U764 ( .A0(n725), .A1(n499), .B0(n674), .Y(n331) );
  AOI2BB2X1 U765 ( .B0(n727), .B1(n468), .A0N(curr_time[16]), .A1N(n688), .Y(
        n680) );
  OAI21XL U766 ( .A0(n724), .A1(n501), .B0(n680), .Y(n323) );
  OAI22XL U767 ( .A0(curr_time[17]), .A1(n683), .B0(n505), .B1(n684), .Y(n682)
         );
  OAI21XL U768 ( .A0(n725), .A1(n525), .B0(n682), .Y(n322) );
  OAI21XL U769 ( .A0(n685), .A1(n684), .B0(curr_time[18]), .Y(n686) );
  OAI22XL U770 ( .A0(curr_time[19]), .A1(n692), .B0(n531), .B1(n693), .Y(n691)
         );
  OAI21XL U771 ( .A0(n725), .A1(n526), .B0(n691), .Y(n320) );
  OAI22XL U772 ( .A0(n724), .A1(n534), .B0(n725), .B1(n510), .Y(n318) );
  OAI22XL U773 ( .A0(n724), .A1(n530), .B0(n725), .B1(n511), .Y(n317) );
  OAI22XL U774 ( .A0(n724), .A1(n502), .B0(n725), .B1(n512), .Y(n316) );
  OAI222XL U775 ( .A0(n696), .A1(n729), .B0(n537), .B1(en_so), .C0(n695), .C1(
        n731), .Y(n338) );
  OAI2BB2XL U776 ( .B0(n696), .B1(n731), .A0N(im_d_w[29]), .A1N(n730), .Y(n337) );
  AOI2BB2X1 U777 ( .B0(\data_path/si_w[9] ), .B1(n727), .A0N(curr_time[9]), 
        .A1N(n708), .Y(n702) );
  OAI21XL U778 ( .A0(n705), .A1(n529), .B0(n702), .Y(n330) );
  OAI2BB2XL U779 ( .B0(n703), .B1(n731), .A0N(im_d_w_9), .A1N(n730), .Y(n357)
         );
  AOI2BB2X1 U780 ( .B0(n466), .B1(n521), .A0N(n466), .A1N(curr_photo_addr[9]), 
        .Y(n400) );
  AOI2BB2X1 U781 ( .B0(n546), .B1(n521), .A0N(n546), .A1N(fb_addr[9]), .Y(n401) );
  OAI21XL U782 ( .A0(curr_time[9]), .A1(n717), .B0(n705), .Y(n706) );
  AOI2BB2X1 U783 ( .B0(n466), .B1(n498), .A0N(n466), .A1N(curr_photo_addr[10]), 
        .Y(n397) );
  AOI2BB2X1 U784 ( .B0(n545), .B1(n498), .A0N(n546), .A1N(fb_addr[10]), .Y(
        n398) );
  AOI2BB1X1 U785 ( .A0N(n711), .A1N(n717), .B0(n726), .Y(n716) );
  AOI2BB2X1 U786 ( .B0(\data_path/si_w[11] ), .B1(n727), .A0N(curr_time[11]), 
        .A1N(n722), .Y(n713) );
  AOI2BB2X1 U787 ( .B0(n466), .B1(n714), .A0N(n466), .A1N(curr_photo_addr[11]), 
        .Y(n394) );
  AOI2BB2X1 U788 ( .B0(n545), .B1(n714), .A0N(n546), .A1N(fb_addr[11]), .Y(
        n395) );
  OAI21XL U789 ( .A0(curr_time[11]), .A1(n717), .B0(n716), .Y(n718) );
  AOI2BB2X1 U790 ( .B0(n466), .B1(n520), .A0N(n466), .A1N(curr_photo_addr[12]), 
        .Y(n391) );
  AOI2BB2X1 U791 ( .B0(n545), .B1(n520), .A0N(en_fb_addr), .A1N(fb_addr[12]), 
        .Y(n392) );
  AOI2BB2X1 U792 ( .B0(n466), .B1(n506), .A0N(n466), .A1N(curr_photo_addr[13]), 
        .Y(n388) );
  AOI2BB2X1 U793 ( .B0(n546), .B1(n506), .A0N(n546), .A1N(fb_addr[13]), .Y(
        n389) );
  AO22X1 U794 ( .A0(\data_path/si_w[13] ), .A1(n734), .B0(n542), .B1(IM_Q[13]), 
        .Y(n390) );
  AO22X1 U795 ( .A0(n727), .A1(\data_path/si_w[14] ), .B0(n726), .B1(
        curr_time[14]), .Y(n325) );
  AOI2BB2X1 U796 ( .B0(n466), .B1(n527), .A0N(n466), .A1N(curr_photo_addr[14]), 
        .Y(n385) );
  AOI2BB2X1 U797 ( .B0(n545), .B1(n527), .A0N(n546), .A1N(fb_addr[14]), .Y(
        n386) );
  AO22X1 U798 ( .A0(\data_path/si_w[14] ), .A1(n734), .B0(n542), .B1(IM_Q[14]), 
        .Y(n387) );
  AO22X1 U799 ( .A0(n727), .A1(\data_path/si_w[15] ), .B0(n726), .B1(
        curr_time[15]), .Y(n324) );
  AOI2BB2X1 U800 ( .B0(n466), .B1(n523), .A0N(n466), .A1N(curr_photo_addr[15]), 
        .Y(n382) );
  AOI2BB2X1 U801 ( .B0(n545), .B1(n523), .A0N(en_fb_addr), .A1N(fb_addr[15]), 
        .Y(n383) );
  AO22X1 U802 ( .A0(\data_path/si_w[15] ), .A1(n734), .B0(n542), .B1(IM_Q[15]), 
        .Y(n384) );
  AOI2BB2X1 U803 ( .B0(n466), .B1(n525), .A0N(n466), .A1N(curr_photo_addr[17]), 
        .Y(n379) );
  AOI2BB2X1 U804 ( .B0(n545), .B1(n525), .A0N(en_fb_addr), .A1N(fb_addr[17]), 
        .Y(n380) );
  AO22X1 U805 ( .A0(\data_path/si_w[17] ), .A1(n734), .B0(n542), .B1(IM_Q[17]), 
        .Y(n381) );
  OAI222XL U806 ( .A0(n732), .A1(n729), .B0(n538), .B1(en_so), .C0(n728), .C1(
        n731), .Y(n348) );
  AOI2BB2X1 U807 ( .B0(n466), .B1(n524), .A0N(n466), .A1N(curr_photo_addr[18]), 
        .Y(n376) );
  AOI2BB2X1 U808 ( .B0(n545), .B1(n524), .A0N(en_fb_addr), .A1N(fb_addr[18]), 
        .Y(n377) );
  AO22X1 U809 ( .A0(\data_path/si_w[18] ), .A1(n734), .B0(n542), .B1(IM_Q[18]), 
        .Y(n378) );
  OAI2BB2XL U810 ( .B0(n732), .B1(n731), .A0N(im_d_w_19), .A1N(n730), .Y(n347)
         );
  AOI2BB2X1 U811 ( .B0(n466), .B1(n526), .A0N(n466), .A1N(curr_photo_addr[19]), 
        .Y(n373) );
  AOI2BB2X1 U812 ( .B0(n545), .B1(n526), .A0N(en_fb_addr), .A1N(fb_addr[19]), 
        .Y(n374) );
  AO22X1 U813 ( .A0(\data_path/si_w[19] ), .A1(n734), .B0(n542), .B1(IM_Q[19]), 
        .Y(n375) );
  AO22X1 U814 ( .A0(\data_path/si_w[20] ), .A1(n734), .B0(n542), .B1(IM_Q[20]), 
        .Y(n372) );
  AO22X1 U815 ( .A0(\data_path/si_w[21] ), .A1(n734), .B0(n542), .B1(IM_Q[21]), 
        .Y(n371) );
  AO22X1 U816 ( .A0(\data_path/si_w[22] ), .A1(n734), .B0(n542), .B1(IM_Q[22]), 
        .Y(n370) );
  AO22X1 U817 ( .A0(\data_path/si_w[23] ), .A1(n734), .B0(n542), .B1(IM_Q[23]), 
        .Y(n369) );
  AO22X1 U818 ( .A0(n466), .A1(n468), .B0(n544), .B1(curr_photo_addr[16]), .Y(
        n11) );
  AO22X1 U819 ( .A0(en_fb_addr), .A1(n468), .B0(n547), .B1(fb_addr[16]), .Y(
        n12) );
  AOI2BB2X1 U820 ( .B0(n466), .B1(n499), .A0N(n466), .A1N(curr_photo_addr[8]), 
        .Y(n13) );
  AOI2BB2X1 U821 ( .B0(n545), .B1(n499), .A0N(n545), .A1N(fb_addr[8]), .Y(n14)
         );
  AOI2BB2X1 U822 ( .B0(n466), .B1(n508), .A0N(n466), .A1N(curr_photo_addr[4]), 
        .Y(n15) );
  AOI2BB2X1 U823 ( .B0(n545), .B1(n508), .A0N(en_fb_addr), .A1N(fb_addr[4]), 
        .Y(n16) );
  AOI2BB2X1 U824 ( .B0(n466), .B1(n509), .A0N(n466), .A1N(curr_photo_addr[2]), 
        .Y(n17) );
  AOI2BB2X1 U825 ( .B0(n545), .B1(n509), .A0N(en_fb_addr), .A1N(fb_addr[2]), 
        .Y(n18) );
  AOI2BB2X1 U826 ( .B0(n466), .B1(n503), .A0N(n466), .A1N(curr_photo_addr[1]), 
        .Y(n19) );
  AOI2BB2X1 U827 ( .B0(n545), .B1(n503), .A0N(en_fb_addr), .A1N(fb_addr[1]), 
        .Y(n20) );
  OAI22XL U828 ( .A0(\data_path/si_w[0] ), .A1(n503), .B0(n514), .B1(
        \data_path/si_w[1] ), .Y(n735) );
  OAI21XL U829 ( .A0(en_curr_photo_size), .A1(n535), .B0(n737), .Y(n23) );
endmodule

