
module CONT ( clk, reset, im_wen_n, cr_a, curr_time, fb_addr, photo_num, 
        curr_photo_addr, curr_photo_size, en_si, en_init_time, en_fb_addr, 
        en_photo_num, en_curr_photo_addr, en_curr_photo_size, en_so, si_sel, 
        init_time_mux_sel, sftr_n, so_mux_sel, expand_sel, \im_a[19]_BAR , 
        \im_a[18]_BAR , \im_a[17]_BAR , \im_a[16]_BAR , \im_a[15]_BAR , 
        \im_a[14]_BAR , \im_a[13]_BAR , \im_a[12]_BAR , \im_a[11]_BAR , 
        \im_a[10]_BAR , \im_a[9]_BAR , \im_a[8]_BAR , \im_a[7]_BAR , 
        \im_a[6]_BAR , \im_a[5]_BAR , \im_a[4]_BAR , \im_a[3]_BAR , 
        \im_a[2]_BAR , \im_a[1]_BAR , \im_a[0]_BAR  );
  output [8:0] cr_a;
  input [23:0] curr_time;
  input [19:0] fb_addr;
  input [1:0] photo_num;
  input [19:0] curr_photo_addr;
  input [1:0] curr_photo_size;
  output [1:0] sftr_n;
  output [1:0] so_mux_sel;
  output [3:0] expand_sel;
  input clk, reset;
  output im_wen_n, en_si, en_init_time, en_fb_addr, en_photo_num,
         en_curr_photo_addr, en_curr_photo_size, en_so, si_sel,
         init_time_mux_sel, \im_a[19]_BAR , \im_a[18]_BAR , \im_a[17]_BAR ,
         \im_a[16]_BAR , \im_a[15]_BAR , \im_a[14]_BAR , \im_a[13]_BAR ,
         \im_a[12]_BAR , \im_a[11]_BAR , \im_a[10]_BAR , \im_a[9]_BAR ,
         \im_a[8]_BAR , \im_a[7]_BAR , \im_a[6]_BAR , \im_a[5]_BAR ,
         \im_a[4]_BAR , \im_a[3]_BAR , \im_a[2]_BAR , \im_a[1]_BAR ,
         \im_a[0]_BAR ;
  wire   n2245, n2246, n2247, n2248, n2249, n2250, \next_write_addr_w[0] ,
         \next_cr_y[0] , \h_0[0] , \m_0[0] , \s_0[0] , N28, N29, N684, N685,
         N686, N687, N688, N689, N690, N691, N910, N911, N912, N913, N914,
         N915, N916, N917, N918, N919, N920, N921, N922, N923, N924, N925,
         N926, N927, N928, N929, N1182, N1183, N1184, N76, next_en_si, N1549,
         N1571, N1591, N1593, \C126/DATA3_0 , \C126/DATA3_1 , \C126/DATA3_2 ,
         \C126/DATA3_3 , \C126/DATA3_4 , \C126/DATA3_5 , \C126/DATA3_6 ,
         \C126/DATA3_7 , \C126/DATA3_8 , \C126/DATA3_9 , \C126/DATA3_10 ,
         \C126/DATA3_11 , \C126/DATA3_12 , \C126/DATA3_13 , \C126/DATA3_14 ,
         \C126/DATA3_15 , \C126/DATA3_16 , \C126/DATA3_17 , \C126/DATA3_18 ,
         n24, n25, n26, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n335, n336,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n351, n352, n353, n354, \DP_OP_436J1_125_1438/n26 ,
         \DP_OP_436J1_125_1438/n25 , \C1/Z_19 , \C1/Z_18 , \C1/Z_17 ,
         \C1/Z_16 , \C1/Z_15 , \C1/Z_14 , \C1/Z_13 , \C1/Z_12 , \C1/Z_11 ,
         \C1/Z_10 , \C1/Z_9 , \C1/Z_8 , \C1/Z_7 , \C1/Z_6 , \C1/Z_5 , \C1/Z_4 ,
         \RSOP_434/C2/CONTROL1 , \C2/Z_18 , \C2/Z_17 , \C2/Z_16 , \C2/Z_15 ,
         \C2/Z_14 , \C2/Z_13 , \C2/Z_12 , \C2/Z_11 , \C2/Z_10 , \C2/Z_9 ,
         \C2/Z_8 , \C2/Z_7 , \C2/Z_6 , \C2/Z_5 , \C2/Z_4 , \C2/Z_3 , \C2/Z_2 ,
         \C2/Z_1 , \C1/Z_3 , \C1/Z_2 , \C1/Z_1 , \C1/Z_0 ,
         \DP_OP_166J1_126_2191/I2 , \DP_OP_166J1_126_2191/I3 ,
         \DP_OP_166J1_126_2191/n27 , \DP_OP_166J1_126_2191/n26 ,
         \DP_OP_166J1_126_2191/n25 , \DP_OP_166J1_126_2191/n24 ,
         \DP_OP_166J1_126_2191/n23 , \DP_OP_166J1_126_2191/n21 ,
         \DP_OP_166J1_126_2191/n17 , \DP_OP_166J1_126_2191/n16 ,
         \DP_OP_166J1_126_2191/n8 , \DP_OP_166J1_126_2191/n7 ,
         \DP_OP_166J1_126_2191/n6 , \DP_OP_166J1_126_2191/n5 ,
         \DP_OP_166J1_126_2191/n4 , \DP_OP_166J1_126_2191/n3 ,
         \DP_OP_166J1_126_2191/n2 , \DP_OP_166J1_126_2191/n1 ,
         \DP_OP_438J1_134_2124/I5 , \DP_OP_438J1_134_2124/n64 ,
         \DP_OP_438J1_134_2124/n63 , \DP_OP_438J1_134_2124/n62 ,
         \DP_OP_438J1_134_2124/n61 , \DP_OP_438J1_134_2124/n60 ,
         \DP_OP_438J1_134_2124/n59 , \DP_OP_438J1_134_2124/n58 ,
         \DP_OP_438J1_134_2124/n57 , \DP_OP_438J1_134_2124/n56 ,
         \DP_OP_438J1_134_2124/n55 , \DP_OP_438J1_134_2124/n54 ,
         \DP_OP_438J1_134_2124/n53 , \DP_OP_438J1_134_2124/n52 ,
         \DP_OP_438J1_134_2124/n51 , \DP_OP_438J1_134_2124/n50 ,
         \DP_OP_438J1_134_2124/n49 , \DP_OP_438J1_134_2124/n48 ,
         \DP_OP_438J1_134_2124/n47 , \DP_OP_438J1_134_2124/n46 ,
         \DP_OP_438J1_134_2124/n40 , \DP_OP_438J1_134_2124/n39 ,
         \DP_OP_438J1_134_2124/n38 , \DP_OP_438J1_134_2124/n37 ,
         \DP_OP_438J1_134_2124/n36 , \DP_OP_438J1_134_2124/n35 ,
         \DP_OP_438J1_134_2124/n34 , \DP_OP_438J1_134_2124/n33 ,
         \DP_OP_438J1_134_2124/n32 , \DP_OP_438J1_134_2124/n31 ,
         \DP_OP_438J1_134_2124/n30 , \DP_OP_438J1_134_2124/n29 ,
         \DP_OP_438J1_134_2124/n28 , \DP_OP_438J1_134_2124/n27 ,
         \DP_OP_438J1_134_2124/n26 , \DP_OP_438J1_134_2124/n25 ,
         \DP_OP_438J1_134_2124/n24 , \DP_OP_438J1_134_2124/n23 ,
         \DP_OP_438J1_134_2124/n22 , \DP_OP_438J1_134_2124/n20 ,
         \DP_OP_438J1_134_2124/n19 , \DP_OP_438J1_134_2124/n18 ,
         \DP_OP_438J1_134_2124/n17 , \DP_OP_438J1_134_2124/n16 ,
         \DP_OP_438J1_134_2124/n15 , \DP_OP_438J1_134_2124/n14 ,
         \DP_OP_438J1_134_2124/n13 , \DP_OP_438J1_134_2124/n12 ,
         \DP_OP_438J1_134_2124/n11 , \DP_OP_438J1_134_2124/n10 ,
         \DP_OP_438J1_134_2124/n9 , \DP_OP_438J1_134_2124/n8 ,
         \DP_OP_438J1_134_2124/n7 , \DP_OP_438J1_134_2124/n6 ,
         \DP_OP_438J1_134_2124/n5 , \DP_OP_438J1_134_2124/n4 ,
         \DP_OP_438J1_134_2124/n3 , \DP_OP_438J1_134_2124/n2 , \intadd_3/A[2] ,
         \intadd_3/A[1] , \intadd_3/A[0] , \intadd_3/B[2] , \intadd_3/B[1] ,
         \intadd_3/B[0] , \intadd_3/CI , \intadd_3/SUM[2] , \intadd_3/SUM[1] ,
         \intadd_3/SUM[0] , \intadd_3/n3 , \intadd_3/n2 , \intadd_3/n1 , n1,
         n2, n3, n4, n5, n6, n8, n10, n12, n14, n16, n18, n20, n22, n27, n29,
         n31, n33, n35, n37, n39, n41, n43, n45, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n147, n148, n149,
         n150, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n184, n186, n188,
         n190, n192, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n337, n338, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244;
  wire   [2:0] next_state;
  wire   [19:0] work_cntr;
  wire   [19:0] next_work_cntr;
  wire   [19:0] global_cntr;
  wire   [19:0] next_glb_cntr;
  wire   [19:0] write_addr;
  wire   [19:0] write_cntr;
  wire   [8:0] next_cr_x;
  wire   [3:0] h_1;
  wire   [3:0] s_1;
  wire   [19:0] read_cntr;
  wire   [8:0] cr_read_cntr;
  wire   [1:0] curr_photo;
  wire   [1:0] next_photo;
  assign \h_0[0]  = curr_time[16];
  assign \m_0[0]  = curr_time[8];
  assign \s_0[0]  = curr_time[0];
  assign en_init_time = N1549;
  assign en_curr_photo_addr = N1571;
  assign en_curr_photo_size = N1591;
  assign init_time_mux_sel = N1593;

  DFFSX1 en_si_reg ( .D(next_en_si), .CK(clk), .SN(n359), .Q(en_si) );
  ADDHXL \DP_OP_166J1_126_2191/U16  ( .A(\C1/Z_0 ), .B(\C1/Z_1 ), .CO(
        \DP_OP_166J1_126_2191/n8 ), .S(\DP_OP_166J1_126_2191/n23 ) );
  ADDFXL \DP_OP_166J1_126_2191/U15  ( .A(\C1/Z_2 ), .B(\C1/Z_1 ), .CI(
        \DP_OP_166J1_126_2191/n8 ), .CO(\DP_OP_166J1_126_2191/n7 ), .S(
        \DP_OP_166J1_126_2191/n24 ) );
  ADDFXL \DP_OP_166J1_126_2191/U14  ( .A(\C1/Z_3 ), .B(\C1/Z_2 ), .CI(
        \DP_OP_166J1_126_2191/n7 ), .CO(\DP_OP_166J1_126_2191/n6 ), .S(
        \DP_OP_166J1_126_2191/n25 ) );
  ADDHXL \DP_OP_166J1_126_2191/U13  ( .A(\C1/Z_3 ), .B(
        \DP_OP_166J1_126_2191/n6 ), .CO(\DP_OP_166J1_126_2191/n27 ), .S(
        \DP_OP_166J1_126_2191/n26 ) );
  AO21X1 \DP_OP_166J1_126_2191/U11  ( .A0(\DP_OP_166J1_126_2191/n23 ), .A1(
        n179), .B0(\DP_OP_166J1_126_2191/I2 ), .Y(\DP_OP_166J1_126_2191/n17 )
         );
  ADDFXL \DP_OP_438J1_134_2124/U61  ( .A(write_addr[1]), .B(fb_addr[1]), .CI(
        \DP_OP_438J1_134_2124/n40 ), .CO(\DP_OP_438J1_134_2124/n39 ), .S(N911)
         );
  ADDFXL \DP_OP_438J1_134_2124/U60  ( .A(write_addr[2]), .B(fb_addr[2]), .CI(
        \DP_OP_438J1_134_2124/n39 ), .CO(\DP_OP_438J1_134_2124/n38 ), .S(N912)
         );
  ADDFXL \DP_OP_438J1_134_2124/U59  ( .A(write_addr[3]), .B(fb_addr[3]), .CI(
        \DP_OP_438J1_134_2124/n38 ), .CO(\DP_OP_438J1_134_2124/n37 ), .S(N913)
         );
  ADDFXL \DP_OP_438J1_134_2124/U58  ( .A(write_addr[4]), .B(fb_addr[4]), .CI(
        \DP_OP_438J1_134_2124/n37 ), .CO(\DP_OP_438J1_134_2124/n36 ), .S(N914)
         );
  ADDFXL \DP_OP_438J1_134_2124/U57  ( .A(write_addr[5]), .B(fb_addr[5]), .CI(
        \DP_OP_438J1_134_2124/n36 ), .CO(\DP_OP_438J1_134_2124/n35 ), .S(N915)
         );
  ADDFXL \DP_OP_438J1_134_2124/U56  ( .A(write_addr[6]), .B(fb_addr[6]), .CI(
        \DP_OP_438J1_134_2124/n35 ), .CO(\DP_OP_438J1_134_2124/n34 ), .S(N916)
         );
  ADDFXL \DP_OP_438J1_134_2124/U55  ( .A(write_addr[7]), .B(fb_addr[7]), .CI(
        \DP_OP_438J1_134_2124/n34 ), .CO(\DP_OP_438J1_134_2124/n33 ), .S(N917)
         );
  ADDFXL \DP_OP_438J1_134_2124/U54  ( .A(n112), .B(fb_addr[8]), .CI(
        \DP_OP_438J1_134_2124/n33 ), .CO(\DP_OP_438J1_134_2124/n32 ), .S(N918)
         );
  ADDFXL \DP_OP_438J1_134_2124/U53  ( .A(n109), .B(fb_addr[9]), .CI(
        \DP_OP_438J1_134_2124/n32 ), .CO(\DP_OP_438J1_134_2124/n31 ), .S(N919)
         );
  ADDFXL \DP_OP_438J1_134_2124/U52  ( .A(n110), .B(fb_addr[10]), .CI(
        \DP_OP_438J1_134_2124/n31 ), .CO(\DP_OP_438J1_134_2124/n30 ), .S(N920)
         );
  ADDFXL \DP_OP_438J1_134_2124/U51  ( .A(write_addr[11]), .B(fb_addr[11]), 
        .CI(\DP_OP_438J1_134_2124/n30 ), .CO(\DP_OP_438J1_134_2124/n29 ), .S(
        N921) );
  ADDFXL \DP_OP_438J1_134_2124/U50  ( .A(write_addr[12]), .B(fb_addr[12]), 
        .CI(\DP_OP_438J1_134_2124/n29 ), .CO(\DP_OP_438J1_134_2124/n28 ), .S(
        N922) );
  ADDFXL \DP_OP_438J1_134_2124/U49  ( .A(write_addr[13]), .B(fb_addr[13]), 
        .CI(\DP_OP_438J1_134_2124/n28 ), .CO(\DP_OP_438J1_134_2124/n27 ), .S(
        N923) );
  ADDFXL \DP_OP_438J1_134_2124/U48  ( .A(write_addr[14]), .B(fb_addr[14]), 
        .CI(\DP_OP_438J1_134_2124/n27 ), .CO(\DP_OP_438J1_134_2124/n26 ), .S(
        N924) );
  ADDFXL \DP_OP_438J1_134_2124/U47  ( .A(write_addr[15]), .B(fb_addr[15]), 
        .CI(\DP_OP_438J1_134_2124/n26 ), .CO(\DP_OP_438J1_134_2124/n25 ), .S(
        N925) );
  ADDFXL \DP_OP_438J1_134_2124/U46  ( .A(write_addr[16]), .B(fb_addr[16]), 
        .CI(\DP_OP_438J1_134_2124/n25 ), .CO(\DP_OP_438J1_134_2124/n24 ), .S(
        N926) );
  ADDFXL \DP_OP_438J1_134_2124/U45  ( .A(write_addr[17]), .B(fb_addr[17]), 
        .CI(\DP_OP_438J1_134_2124/n24 ), .CO(\DP_OP_438J1_134_2124/n23 ), .S(
        N927) );
  ADDFXL \DP_OP_438J1_134_2124/U44  ( .A(write_addr[18]), .B(fb_addr[18]), 
        .CI(\DP_OP_438J1_134_2124/n23 ), .CO(\DP_OP_438J1_134_2124/n22 ), .S(
        N928) );
  AO22X1 \DP_OP_438J1_134_2124/U40  ( .A0(N911), .A1(si_sel), .B0(
        \DP_OP_438J1_134_2124/I5 ), .B1(\C2/Z_1 ), .Y(
        \DP_OP_438J1_134_2124/n46 ) );
  AO22X1 \DP_OP_438J1_134_2124/U39  ( .A0(N912), .A1(si_sel), .B0(
        \DP_OP_438J1_134_2124/I5 ), .B1(\C2/Z_2 ), .Y(
        \DP_OP_438J1_134_2124/n47 ) );
  AO22X1 \DP_OP_438J1_134_2124/U38  ( .A0(N913), .A1(si_sel), .B0(
        \DP_OP_438J1_134_2124/I5 ), .B1(\C2/Z_3 ), .Y(
        \DP_OP_438J1_134_2124/n48 ) );
  AO22X1 \DP_OP_438J1_134_2124/U37  ( .A0(N914), .A1(si_sel), .B0(
        \DP_OP_438J1_134_2124/I5 ), .B1(\C2/Z_4 ), .Y(
        \DP_OP_438J1_134_2124/n49 ) );
  AO22X1 \DP_OP_438J1_134_2124/U36  ( .A0(N915), .A1(si_sel), .B0(
        \DP_OP_438J1_134_2124/I5 ), .B1(\C2/Z_5 ), .Y(
        \DP_OP_438J1_134_2124/n50 ) );
  AO22X1 \DP_OP_438J1_134_2124/U35  ( .A0(N916), .A1(si_sel), .B0(
        \DP_OP_438J1_134_2124/I5 ), .B1(\C2/Z_6 ), .Y(
        \DP_OP_438J1_134_2124/n51 ) );
  AO22X1 \DP_OP_438J1_134_2124/U34  ( .A0(N917), .A1(si_sel), .B0(
        \DP_OP_438J1_134_2124/I5 ), .B1(\C2/Z_7 ), .Y(
        \DP_OP_438J1_134_2124/n52 ) );
  AO22X1 \DP_OP_438J1_134_2124/U33  ( .A0(N918), .A1(si_sel), .B0(
        \DP_OP_438J1_134_2124/I5 ), .B1(\C2/Z_8 ), .Y(
        \DP_OP_438J1_134_2124/n53 ) );
  AO22X1 \DP_OP_438J1_134_2124/U32  ( .A0(N919), .A1(si_sel), .B0(
        \DP_OP_438J1_134_2124/I5 ), .B1(\C2/Z_9 ), .Y(
        \DP_OP_438J1_134_2124/n54 ) );
  AO22X1 \DP_OP_438J1_134_2124/U31  ( .A0(N920), .A1(si_sel), .B0(
        \DP_OP_438J1_134_2124/I5 ), .B1(\C2/Z_10 ), .Y(
        \DP_OP_438J1_134_2124/n55 ) );
  AO22X1 \DP_OP_438J1_134_2124/U30  ( .A0(N921), .A1(si_sel), .B0(
        \DP_OP_438J1_134_2124/I5 ), .B1(\C2/Z_11 ), .Y(
        \DP_OP_438J1_134_2124/n56 ) );
  AO22X1 \DP_OP_438J1_134_2124/U29  ( .A0(N922), .A1(si_sel), .B0(
        \DP_OP_438J1_134_2124/I5 ), .B1(\C2/Z_12 ), .Y(
        \DP_OP_438J1_134_2124/n57 ) );
  AO22X1 \DP_OP_438J1_134_2124/U28  ( .A0(N923), .A1(si_sel), .B0(
        \DP_OP_438J1_134_2124/I5 ), .B1(\C2/Z_13 ), .Y(
        \DP_OP_438J1_134_2124/n58 ) );
  AO22X1 \DP_OP_438J1_134_2124/U27  ( .A0(N924), .A1(si_sel), .B0(
        \DP_OP_438J1_134_2124/I5 ), .B1(\C2/Z_14 ), .Y(
        \DP_OP_438J1_134_2124/n59 ) );
  AO22X1 \DP_OP_438J1_134_2124/U26  ( .A0(N925), .A1(si_sel), .B0(
        \DP_OP_438J1_134_2124/I5 ), .B1(\C2/Z_15 ), .Y(
        \DP_OP_438J1_134_2124/n60 ) );
  AO22X1 \DP_OP_438J1_134_2124/U25  ( .A0(N926), .A1(si_sel), .B0(
        \DP_OP_438J1_134_2124/I5 ), .B1(\C2/Z_16 ), .Y(
        \DP_OP_438J1_134_2124/n61 ) );
  AO22X1 \DP_OP_438J1_134_2124/U24  ( .A0(N927), .A1(si_sel), .B0(
        \DP_OP_438J1_134_2124/I5 ), .B1(\C2/Z_17 ), .Y(
        \DP_OP_438J1_134_2124/n62 ) );
  AO22X1 \DP_OP_438J1_134_2124/U23  ( .A0(N928), .A1(si_sel), .B0(
        \DP_OP_438J1_134_2124/I5 ), .B1(\C2/Z_18 ), .Y(
        \DP_OP_438J1_134_2124/n63 ) );
  ADDFXL \DP_OP_438J1_134_2124/U20  ( .A(\DP_OP_438J1_134_2124/n20 ), .B(n627), 
        .CI(\DP_OP_438J1_134_2124/n46 ), .CO(\DP_OP_438J1_134_2124/n19 ), .S(
        \C126/DATA3_1 ) );
  ADDFXL \DP_OP_438J1_134_2124/U19  ( .A(\DP_OP_438J1_134_2124/n47 ), .B(n628), 
        .CI(\DP_OP_438J1_134_2124/n19 ), .CO(\DP_OP_438J1_134_2124/n18 ), .S(
        \C126/DATA3_2 ) );
  ADDFXL \DP_OP_438J1_134_2124/U18  ( .A(\DP_OP_438J1_134_2124/n48 ), .B(n629), 
        .CI(\DP_OP_438J1_134_2124/n18 ), .CO(\DP_OP_438J1_134_2124/n17 ), .S(
        \C126/DATA3_3 ) );
  ADDFXL \DP_OP_438J1_134_2124/U17  ( .A(\DP_OP_438J1_134_2124/n49 ), .B(
        \C1/Z_4 ), .CI(\DP_OP_438J1_134_2124/n17 ), .CO(
        \DP_OP_438J1_134_2124/n16 ), .S(\C126/DATA3_4 ) );
  ADDFXL \DP_OP_438J1_134_2124/U16  ( .A(\DP_OP_438J1_134_2124/n50 ), .B(
        \C1/Z_5 ), .CI(\DP_OP_438J1_134_2124/n16 ), .CO(
        \DP_OP_438J1_134_2124/n15 ), .S(\C126/DATA3_5 ) );
  ADDFXL \DP_OP_438J1_134_2124/U15  ( .A(\DP_OP_438J1_134_2124/n51 ), .B(
        \C1/Z_6 ), .CI(\DP_OP_438J1_134_2124/n15 ), .CO(
        \DP_OP_438J1_134_2124/n14 ), .S(\C126/DATA3_6 ) );
  ADDFXL \DP_OP_438J1_134_2124/U14  ( .A(\DP_OP_438J1_134_2124/n52 ), .B(
        \C1/Z_7 ), .CI(\DP_OP_438J1_134_2124/n14 ), .CO(
        \DP_OP_438J1_134_2124/n13 ), .S(\C126/DATA3_7 ) );
  ADDFXL \DP_OP_438J1_134_2124/U13  ( .A(\DP_OP_438J1_134_2124/n53 ), .B(
        \C1/Z_8 ), .CI(\DP_OP_438J1_134_2124/n13 ), .CO(
        \DP_OP_438J1_134_2124/n12 ), .S(\C126/DATA3_8 ) );
  ADDFXL \DP_OP_438J1_134_2124/U12  ( .A(\DP_OP_438J1_134_2124/n54 ), .B(
        \C1/Z_9 ), .CI(\DP_OP_438J1_134_2124/n12 ), .CO(
        \DP_OP_438J1_134_2124/n11 ), .S(\C126/DATA3_9 ) );
  ADDFXL \DP_OP_438J1_134_2124/U11  ( .A(\DP_OP_438J1_134_2124/n55 ), .B(
        \C1/Z_10 ), .CI(\DP_OP_438J1_134_2124/n11 ), .CO(
        \DP_OP_438J1_134_2124/n10 ), .S(\C126/DATA3_10 ) );
  ADDFXL \DP_OP_438J1_134_2124/U10  ( .A(\DP_OP_438J1_134_2124/n56 ), .B(
        \C1/Z_11 ), .CI(\DP_OP_438J1_134_2124/n10 ), .CO(
        \DP_OP_438J1_134_2124/n9 ), .S(\C126/DATA3_11 ) );
  ADDFXL \DP_OP_438J1_134_2124/U9  ( .A(\DP_OP_438J1_134_2124/n57 ), .B(
        \C1/Z_12 ), .CI(\DP_OP_438J1_134_2124/n9 ), .CO(
        \DP_OP_438J1_134_2124/n8 ), .S(\C126/DATA3_12 ) );
  ADDFXL \DP_OP_438J1_134_2124/U8  ( .A(\DP_OP_438J1_134_2124/n58 ), .B(
        \C1/Z_13 ), .CI(\DP_OP_438J1_134_2124/n8 ), .CO(
        \DP_OP_438J1_134_2124/n7 ), .S(\C126/DATA3_13 ) );
  ADDFXL \DP_OP_438J1_134_2124/U7  ( .A(\DP_OP_438J1_134_2124/n59 ), .B(
        \C1/Z_14 ), .CI(\DP_OP_438J1_134_2124/n7 ), .CO(
        \DP_OP_438J1_134_2124/n6 ), .S(\C126/DATA3_14 ) );
  ADDFXL \DP_OP_438J1_134_2124/U6  ( .A(\DP_OP_438J1_134_2124/n60 ), .B(
        \C1/Z_15 ), .CI(\DP_OP_438J1_134_2124/n6 ), .CO(
        \DP_OP_438J1_134_2124/n5 ), .S(\C126/DATA3_15 ) );
  ADDFXL \DP_OP_438J1_134_2124/U5  ( .A(\DP_OP_438J1_134_2124/n61 ), .B(
        \C1/Z_16 ), .CI(\DP_OP_438J1_134_2124/n5 ), .CO(
        \DP_OP_438J1_134_2124/n4 ), .S(\C126/DATA3_16 ) );
  ADDFXL \DP_OP_438J1_134_2124/U4  ( .A(\DP_OP_438J1_134_2124/n62 ), .B(
        \C1/Z_17 ), .CI(\DP_OP_438J1_134_2124/n4 ), .CO(
        \DP_OP_438J1_134_2124/n3 ), .S(\C126/DATA3_17 ) );
  ADDFXL \DP_OP_438J1_134_2124/U3  ( .A(\DP_OP_438J1_134_2124/n63 ), .B(
        \C1/Z_18 ), .CI(\DP_OP_438J1_134_2124/n3 ), .CO(
        \DP_OP_438J1_134_2124/n2 ), .S(\C126/DATA3_18 ) );
  ADDFXL \intadd_3/U4  ( .A(\intadd_3/A[0] ), .B(\intadd_3/B[0] ), .CI(
        \intadd_3/CI ), .CO(\intadd_3/n3 ), .S(\intadd_3/SUM[0] ) );
  ADDFXL \intadd_3/U3  ( .A(\intadd_3/A[1] ), .B(\intadd_3/B[1] ), .CI(
        \intadd_3/n3 ), .CO(\intadd_3/n2 ), .S(\intadd_3/SUM[1] ) );
  DFFRX1 \write_addr_reg/q_reg[0]  ( .D(n307), .CK(clk), .RN(n357), .Q(
        \next_write_addr_w[0] ), .QN(n330) );
  DFFRX1 \cr_read_cntr_reg/q_reg[1]  ( .D(n315), .CK(clk), .RN(n358), .Q(N685), 
        .QN(n323) );
  DFFRX1 \cr_read_cntr_reg/q_reg[7]  ( .D(n309), .CK(clk), .RN(n358), .Q(
        cr_read_cntr[7]), .QN(n287) );
  DFFRX1 \cr_read_cntr_reg/q_reg[6]  ( .D(n310), .CK(clk), .RN(n358), .Q(
        cr_read_cntr[6]), .QN(n286) );
  DFFRX1 \write_addr_reg/q_reg[12]  ( .D(n295), .CK(clk), .RN(n357), .Q(
        write_addr[12]), .QN(n275) );
  DFFRX1 \cr_read_cntr_reg/q_reg[3]  ( .D(n313), .CK(clk), .RN(n358), .Q(
        cr_read_cntr[3]), .QN(n240) );
  DFFRX1 \write_addr_reg/q_reg[5]  ( .D(n302), .CK(clk), .RN(n358), .Q(
        write_addr[5]), .QN(n239) );
  DFFRX1 \write_addr_reg/q_reg[3]  ( .D(n304), .CK(clk), .RN(n358), .Q(
        write_addr[3]), .QN(n238) );
  DFFRX1 \cr_read_cntr_reg/q_reg[2]  ( .D(n314), .CK(clk), .RN(n358), .Q(N686), 
        .QN(n224) );
  DFFRX1 \read_cntr_reg/q_reg[0]  ( .D(n336), .CK(clk), .RN(n358), .Q(
        read_cntr[0]), .QN(n277) );
  DFFRX1 \read_cntr_reg/q_reg[1]  ( .D(n335), .CK(clk), .RN(n357), .Q(
        read_cntr[1]), .QN(n326) );
  DFFRX1 \write_addr_reg/q_reg[7]  ( .D(n300), .CK(clk), .RN(n357), .Q(
        write_addr[7]), .QN(n328) );
  DFFRX1 \write_addr_reg/q_reg[4]  ( .D(n303), .CK(clk), .RN(n114), .Q(
        write_addr[4]), .QN(n281) );
  DFFRX1 \write_addr_reg/q_reg[2]  ( .D(n305), .CK(clk), .RN(n357), .Q(
        write_addr[2]), .QN(n329) );
  DFFRX1 \state_reg[1]  ( .D(next_state[1]), .CK(clk), .RN(n357), .QN(n25) );
  ADDHXL \DP_OP_166J1_126_2191/U6  ( .A(N28), .B(\DP_OP_166J1_126_2191/n16 ), 
        .CO(\DP_OP_166J1_126_2191/n5 ), .S(N687) );
  AND2XL \DP_OP_166J1_126_2191/U12  ( .A(\C1/Z_0 ), .B(n179), .Y(
        \DP_OP_166J1_126_2191/n16 ) );
  AND2XL \DP_OP_166J1_126_2191/U7  ( .A(\DP_OP_166J1_126_2191/n27 ), .B(n179), 
        .Y(\DP_OP_166J1_126_2191/n21 ) );
  DFFSX2 \state_reg[0]  ( .D(n635), .CK(clk), .SN(n359), .Q(n26), .QN(n252) );
  ADDFX2 \intadd_3/U2  ( .A(\intadd_3/A[2] ), .B(\intadd_3/B[2] ), .CI(
        \intadd_3/n2 ), .CO(\intadd_3/n1 ), .S(\intadd_3/SUM[2] ) );
  ADDHX1 \DP_OP_438J1_134_2124/U62  ( .A(fb_addr[0]), .B(
        \next_write_addr_w[0] ), .CO(\DP_OP_438J1_134_2124/n40 ), .S(N910) );
  DFFRX1 \global_cntr_reg[8]  ( .D(n650), .CK(clk), .RN(n114), .Q(
        global_cntr[8]), .QN(n579) );
  DFFRX1 \global_cntr_reg[19]  ( .D(n638), .CK(clk), .RN(n359), .Q(
        global_cntr[19]) );
  DFFRX1 \write_cntr_reg/q_reg[2]  ( .D(n353), .CK(clk), .RN(n114), .Q(
        write_cntr[2]) );
  DFFRX1 \write_addr_reg/q_reg[15]  ( .D(n292), .CK(clk), .RN(n358), .Q(
        write_addr[15]), .QN(n2203) );
  DFFRX1 \cr_read_cntr_reg/q_reg[5]  ( .D(n311), .CK(clk), .RN(n114), .Q(
        cr_read_cntr[5]) );
  DFFRX1 \cr_read_cntr_reg/q_reg[8]  ( .D(n308), .CK(clk), .RN(n357), .Q(
        cr_read_cntr[8]) );
  DFFRX1 \global_cntr_reg[0]  ( .D(n279), .CK(clk), .RN(n359), .Q(
        global_cntr[0]), .QN(n279) );
  DFFRX1 \global_cntr_reg[2]  ( .D(next_glb_cntr[2]), .CK(clk), .RN(n359), .Q(
        global_cntr[2]), .QN(n226) );
  DFFRX1 \write_cntr_reg/q_reg[10]  ( .D(n343), .CK(clk), .RN(n358), .Q(
        write_cntr[10]), .QN(n221) );
  DFFRX1 \write_cntr_reg/q_reg[7]  ( .D(n345), .CK(clk), .RN(n114), .Q(
        write_cntr[7]), .QN(n256) );
  DFFRX1 \cr_read_cntr_reg/q_reg[4]  ( .D(n312), .CK(clk), .RN(n114), .Q(
        cr_read_cntr[4]), .QN(n322) );
  DFFSRX1 \global_cntr_reg[3]  ( .D(n655), .CK(clk), .SN(1'b1), .RN(n357), .Q(
        global_cntr[3]), .QN(n280) );
  DFFSRX1 \global_cntr_reg[4]  ( .D(n654), .CK(clk), .SN(1'b1), .RN(n114), .Q(
        global_cntr[4]), .QN(n282) );
  DFFSRX1 \global_cntr_reg[5]  ( .D(n653), .CK(clk), .SN(1'b1), .RN(n358), .Q(
        global_cntr[5]), .QN(n241) );
  DFFSRX1 \global_cntr_reg[6]  ( .D(next_glb_cntr[6]), .CK(clk), .SN(1'b1), 
        .RN(n114), .Q(global_cntr[6]), .QN(n246) );
  DFFSRX1 \global_cntr_reg[7]  ( .D(n651), .CK(clk), .SN(1'b1), .RN(n357), .Q(
        global_cntr[7]), .QN(n283) );
  DFFSRX1 \global_cntr_reg[9]  ( .D(n649), .CK(clk), .SN(1'b1), .RN(n114), .Q(
        global_cntr[9]), .QN(n233) );
  DFFSRX1 \global_cntr_reg[10]  ( .D(n647), .CK(clk), .SN(1'b1), .RN(n358), 
        .Q(global_cntr[10]), .QN(n284) );
  DFFSRX1 \global_cntr_reg[11]  ( .D(n646), .CK(clk), .SN(1'b1), .RN(n114), 
        .Q(global_cntr[11]), .QN(n250) );
  DFFSRX1 \global_cntr_reg[12]  ( .D(n645), .CK(clk), .SN(1'b1), .RN(n357), 
        .Q(global_cntr[12]), .QN(n244) );
  DFFSRX1 \global_cntr_reg[13]  ( .D(n644), .CK(clk), .SN(1'b1), .RN(n114), 
        .Q(global_cntr[13]), .QN(n317) );
  DFFSRX1 \global_cntr_reg[14]  ( .D(n643), .CK(clk), .SN(1'b1), .RN(n358), 
        .Q(global_cntr[14]), .QN(n243) );
  DFFSRX1 \global_cntr_reg[15]  ( .D(n642), .CK(clk), .SN(1'b1), .RN(n114), 
        .Q(global_cntr[15]), .QN(n319) );
  DFFSRX1 \global_cntr_reg[16]  ( .D(n641), .CK(clk), .SN(1'b1), .RN(n357), 
        .Q(global_cntr[16]), .QN(n225) );
  DFFSRX1 \global_cntr_reg[18]  ( .D(n639), .CK(clk), .SN(1'b1), .RN(n114), 
        .Q(global_cntr[18]), .QN(n247) );
  DFFSRX1 \state_reg[2]  ( .D(next_state[2]), .CK(clk), .SN(1'b1), .RN(n358), 
        .Q(n234), .QN(n24) );
  DFFSRX1 \curr_photo_reg[1]  ( .D(next_photo[1]), .CK(clk), .SN(1'b1), .RN(
        n114), .Q(curr_photo[1]), .QN(n325) );
  DFFSRX1 \curr_photo_reg[0]  ( .D(next_photo[0]), .CK(clk), .SN(1'b1), .RN(
        n357), .Q(curr_photo[0]), .QN(n331) );
  DFFSRX1 \write_addr_reg/q_reg[18]  ( .D(n289), .CK(clk), .SN(1'b1), .RN(n114), .Q(write_addr[18]), .QN(n321) );
  DFFSRX1 \write_cntr_reg/q_reg[0]  ( .D(n349), .CK(clk), .SN(1'b1), .RN(n358), 
        .Q(write_cntr[0]), .QN(n272) );
  DFFSRX1 \write_cntr_reg/q_reg[14]  ( .D(n339), .CK(clk), .SN(1'b1), .RN(n114), .Q(write_cntr[14]), .QN(n254) );
  DFFSRX1 \write_cntr_reg/q_reg[11]  ( .D(n342), .CK(clk), .SN(1'b1), .RN(n357), .Q(write_cntr[11]), .QN(n248) );
  DFFSRX1 \write_cntr_reg/q_reg[9]  ( .D(n344), .CK(clk), .SN(1'b1), .RN(n114), 
        .Q(write_cntr[9]), .QN(n230) );
  DFFSRX1 \write_cntr_reg/q_reg[4]  ( .D(n352), .CK(clk), .SN(1'b1), .RN(n358), 
        .Q(write_cntr[4]), .QN(n285) );
  DFFSRX1 \write_addr_reg/q_reg[19]  ( .D(n288), .CK(clk), .SN(1'b1), .RN(n114), .Q(write_addr[19]), .QN(n276) );
  DFFSRX1 \write_addr_reg/q_reg[17]  ( .D(n290), .CK(clk), .SN(1'b1), .RN(n357), .Q(write_addr[17]), .QN(n318) );
  DFFSRX1 \write_addr_reg/q_reg[14]  ( .D(n293), .CK(clk), .SN(1'b1), .RN(n114), .Q(write_addr[14]), .QN(n274) );
  DFFSRX1 \write_cntr_reg/q_reg[1]  ( .D(n354), .CK(clk), .SN(1'b1), .RN(n358), 
        .Q(write_cntr[1]), .QN(n271) );
  DFFSRX1 \write_cntr_reg/q_reg[13]  ( .D(n340), .CK(clk), .SN(1'b1), .RN(n114), .Q(write_cntr[13]), .QN(n324) );
  DFFSRX1 \write_cntr_reg/q_reg[3]  ( .D(n348), .CK(clk), .SN(1'b1), .RN(n357), 
        .Q(write_cntr[3]), .QN(n270) );
  DFFSRX1 \write_cntr_reg/q_reg[8]  ( .D(n351), .CK(clk), .SN(1'b1), .RN(n114), 
        .Q(write_cntr[8]), .QN(n245) );
  DFFSRX1 \write_cntr_reg/q_reg[5]  ( .D(n347), .CK(clk), .SN(1'b1), .RN(n358), 
        .Q(write_cntr[5]), .QN(n253) );
  DFFSRX1 \cr_read_cntr_reg/q_reg[0]  ( .D(n316), .CK(clk), .SN(1'b1), .RN(
        n114), .Q(N684), .QN(n231) );
  DFFRX2 \write_cntr_reg/q_reg[6]  ( .D(n346), .CK(clk), .RN(n358), .Q(
        write_cntr[6]) );
  DFFRX2 \write_addr_reg/q_reg[1]  ( .D(n306), .CK(clk), .RN(n358), .Q(
        write_addr[1]) );
  DFFRX2 \write_addr_reg/q_reg[6]  ( .D(n301), .CK(clk), .RN(n358), .Q(
        write_addr[6]) );
  DFFRX2 \write_addr_reg/q_reg[11]  ( .D(n296), .CK(clk), .RN(n358), .Q(
        write_addr[11]) );
  DFFRX2 \write_addr_reg/q_reg[13]  ( .D(n294), .CK(clk), .RN(n359), .Q(
        write_addr[13]) );
  DFFRX4 \work_cntr_reg[2]  ( .D(next_work_cntr[2]), .CK(clk), .RN(n357), .Q(
        N1183), .QN(n257) );
  DFFRX4 \work_cntr_reg[6]  ( .D(next_work_cntr[6]), .CK(clk), .RN(n359), .Q(
        work_cntr[6]), .QN(n263) );
  DFFRX4 \work_cntr_reg[4]  ( .D(next_work_cntr[4]), .CK(clk), .RN(n114), .Q(
        work_cntr[4]), .QN(n223) );
  DFFRX4 \work_cntr_reg[15]  ( .D(next_work_cntr[15]), .CK(clk), .RN(n357), 
        .Q(work_cntr[15]), .QN(n264) );
  DFFRX2 \work_cntr_reg[0]  ( .D(n153), .CK(clk), .RN(n357), .Q(N76), .QN(n258) );
  DFFRX2 \work_cntr_reg[9]  ( .D(next_work_cntr[9]), .CK(clk), .RN(n359), .Q(
        work_cntr[9]), .QN(n265) );
  DFFRX2 \work_cntr_reg[12]  ( .D(next_work_cntr[12]), .CK(clk), .RN(n114), 
        .Q(work_cntr[12]), .QN(n209) );
  DFFRX2 \work_cntr_reg[7]  ( .D(next_work_cntr[7]), .CK(clk), .RN(n114), .Q(
        work_cntr[7]), .QN(n261) );
  DFFRX2 \work_cntr_reg[10]  ( .D(next_work_cntr[10]), .CK(clk), .RN(n357), 
        .Q(work_cntr[10]), .QN(n269) );
  DFFRX2 \work_cntr_reg[11]  ( .D(next_work_cntr[11]), .CK(clk), .RN(n359), 
        .Q(work_cntr[11]), .QN(n267) );
  DFFRX2 \work_cntr_reg[16]  ( .D(next_work_cntr[16]), .CK(clk), .RN(n357), 
        .Q(work_cntr[16]), .QN(n260) );
  DFFRX2 \work_cntr_reg[17]  ( .D(next_work_cntr[17]), .CK(clk), .RN(n114), 
        .Q(work_cntr[17]), .QN(n222) );
  DFFRX2 \work_cntr_reg[13]  ( .D(next_work_cntr[13]), .CK(clk), .RN(n359), 
        .Q(work_cntr[13]), .QN(n268) );
  DFFRX2 \work_cntr_reg[3]  ( .D(next_work_cntr[3]), .CK(clk), .RN(n114), .Q(
        N1184), .QN(n228) );
  DFFRX2 \work_cntr_reg[19]  ( .D(next_work_cntr[19]), .CK(clk), .RN(n114), 
        .Q(work_cntr[19]), .QN(n259) );
  DFFRX2 \work_cntr_reg[18]  ( .D(next_work_cntr[18]), .CK(clk), .RN(n114), 
        .Q(work_cntr[18]), .QN(n236) );
  DFFRX2 \work_cntr_reg[5]  ( .D(next_work_cntr[5]), .CK(clk), .RN(n114), .Q(
        work_cntr[5]), .QN(n229) );
  DFFRXL \write_addr_reg/q_reg[8]  ( .D(n299), .CK(clk), .RN(n358), .Q(
        write_addr[8]), .QN(n278) );
  DFFRX2 \write_cntr_reg/q_reg[12]  ( .D(n341), .CK(clk), .RN(n114), .Q(
        write_cntr[12]), .QN(n235) );
  DFFRX2 \global_cntr_reg[1]  ( .D(next_glb_cntr[1]), .CK(clk), .RN(n114), .Q(
        global_cntr[1]), .QN(n249) );
  DFFRX2 \work_cntr_reg[8]  ( .D(next_work_cntr[8]), .CK(clk), .RN(n114), .Q(
        work_cntr[8]), .QN(n262) );
  DFFRXL \write_addr_reg/q_reg[10]  ( .D(n297), .CK(clk), .RN(n114), .Q(
        write_addr[10]), .QN(n327) );
  DFFRXL \write_addr_reg/q_reg[9]  ( .D(n298), .CK(clk), .RN(n357), .Q(
        write_addr[9]), .QN(n273) );
  DFFRXL \global_cntr_reg[17]  ( .D(n640), .CK(clk), .RN(n114), .Q(
        global_cntr[17]), .QN(n320) );
  DFFRX1 \work_cntr_reg[14]  ( .D(next_work_cntr[14]), .CK(clk), .RN(n359), 
        .Q(work_cntr[14]) );
  DFFRX1 \write_addr_reg/q_reg[16]  ( .D(n291), .CK(clk), .RN(n359), .Q(
        write_addr[16]), .QN(n2230) );
  DFFRX2 \work_cntr_reg[1]  ( .D(next_work_cntr[1]), .CK(clk), .RN(n357), .Q(
        N1182), .QN(n227) );
  ADDFX2 \DP_OP_166J1_126_2191/U5  ( .A(\DP_OP_166J1_126_2191/n5 ), .B(N29), 
        .CI(\DP_OP_166J1_126_2191/n17 ), .CO(\DP_OP_166J1_126_2191/n4 ), .S(
        N688) );
  AND2X2 U3 ( .A(n478), .B(n485), .Y(n1) );
  OR2X1 U4 ( .A(n1534), .B(n1535), .Y(n196) );
  AOI2BB2X1 U5 ( .B0(n1978), .B1(n2152), .A0N(n1978), .A1N(n2152), .Y(n786) );
  AOI2BB2X1 U6 ( .B0(n1447), .B1(n713), .A0N(n1447), .A1N(n713), .Y(n903) );
  AOI2BB2X1 U7 ( .B0(n908), .B1(n907), .A0N(n908), .A1N(n907), .Y(n1980) );
  OA22X1 U8 ( .A0(n1), .A1(n479), .B0(n480), .B1(n484), .Y(n512) );
  NAND2X1 U9 ( .A(n1277), .B(n1438), .Y(n1440) );
  AND2X2 U10 ( .A(im_wen_n), .B(n220), .Y(n266) );
  BUFX4 U11 ( .A(n266), .Y(n147) );
  NAND2X4 U12 ( .A(en_so), .B(n252), .Y(n2241) );
  OR2X1 U13 ( .A(n231), .B(n2241), .Y(n2) );
  OR2X1 U14 ( .A(n323), .B(n2241), .Y(n3) );
  OR2X1 U15 ( .A(n224), .B(n2241), .Y(n4) );
  OR2X1 U16 ( .A(n6), .B(n2241), .Y(n5) );
  XNOR2X1 U17 ( .A(\DP_OP_166J1_126_2191/n1 ), .B(\DP_OP_166J1_126_2191/n21 ), 
        .Y(n6) );
  AOI21X1 U18 ( .A0(n626), .A1(\C126/DATA3_0 ), .B0(n8), .Y(\im_a[0]_BAR ) );
  AO22X1 U19 ( .A0(n356), .A1(N910), .B0(n337), .B1(global_cntr[0]), .Y(n8) );
  AOI21X1 U20 ( .A0(n626), .A1(\C126/DATA3_1 ), .B0(n10), .Y(\im_a[1]_BAR ) );
  AO22X1 U21 ( .A0(n356), .A1(N911), .B0(n337), .B1(global_cntr[1]), .Y(n10)
         );
  AOI21X1 U22 ( .A0(n626), .A1(\C126/DATA3_2 ), .B0(n12), .Y(\im_a[2]_BAR ) );
  AO22X1 U23 ( .A0(n625), .A1(N912), .B0(n337), .B1(global_cntr[2]), .Y(n12)
         );
  AOI21X1 U24 ( .A0(n626), .A1(\C126/DATA3_3 ), .B0(n14), .Y(\im_a[3]_BAR ) );
  AO22X1 U25 ( .A0(n356), .A1(N913), .B0(n337), .B1(global_cntr[3]), .Y(n14)
         );
  AOI21X1 U26 ( .A0(n626), .A1(\C126/DATA3_4 ), .B0(n16), .Y(\im_a[4]_BAR ) );
  AO22X1 U27 ( .A0(n356), .A1(N914), .B0(n337), .B1(global_cntr[4]), .Y(n16)
         );
  AOI21X1 U28 ( .A0(n626), .A1(\C126/DATA3_5 ), .B0(n18), .Y(\im_a[5]_BAR ) );
  AO22X1 U29 ( .A0(n625), .A1(N915), .B0(n337), .B1(global_cntr[5]), .Y(n18)
         );
  AOI21X1 U30 ( .A0(n626), .A1(\C126/DATA3_6 ), .B0(n20), .Y(\im_a[6]_BAR ) );
  AO22X1 U31 ( .A0(n625), .A1(N916), .B0(n337), .B1(global_cntr[6]), .Y(n20)
         );
  AOI21X1 U32 ( .A0(n626), .A1(\C126/DATA3_7 ), .B0(n22), .Y(\im_a[7]_BAR ) );
  AO22X1 U33 ( .A0(n356), .A1(N917), .B0(n337), .B1(global_cntr[7]), .Y(n22)
         );
  AOI21X1 U34 ( .A0(n626), .A1(\C126/DATA3_8 ), .B0(n27), .Y(\im_a[8]_BAR ) );
  AO22X1 U35 ( .A0(n356), .A1(N918), .B0(n337), .B1(global_cntr[8]), .Y(n27)
         );
  AOI21X1 U36 ( .A0(n626), .A1(\C126/DATA3_9 ), .B0(n29), .Y(\im_a[9]_BAR ) );
  AO22X1 U37 ( .A0(n356), .A1(N919), .B0(n337), .B1(global_cntr[9]), .Y(n29)
         );
  AOI21X1 U38 ( .A0(n626), .A1(\C126/DATA3_10 ), .B0(n31), .Y(\im_a[10]_BAR )
         );
  AO22X1 U39 ( .A0(n625), .A1(N920), .B0(n337), .B1(global_cntr[10]), .Y(n31)
         );
  AOI21X1 U40 ( .A0(n626), .A1(\C126/DATA3_11 ), .B0(n33), .Y(\im_a[11]_BAR )
         );
  AO22X1 U41 ( .A0(n356), .A1(N921), .B0(n337), .B1(global_cntr[11]), .Y(n33)
         );
  AOI21X1 U42 ( .A0(n626), .A1(\C126/DATA3_12 ), .B0(n35), .Y(\im_a[12]_BAR )
         );
  AO22X1 U43 ( .A0(n356), .A1(N922), .B0(n337), .B1(global_cntr[12]), .Y(n35)
         );
  AOI21X1 U44 ( .A0(n626), .A1(\C126/DATA3_13 ), .B0(n37), .Y(\im_a[13]_BAR )
         );
  AO22X1 U45 ( .A0(n356), .A1(N923), .B0(n337), .B1(global_cntr[13]), .Y(n37)
         );
  AOI21X1 U46 ( .A0(n626), .A1(\C126/DATA3_14 ), .B0(n39), .Y(\im_a[14]_BAR )
         );
  AO22X1 U47 ( .A0(n625), .A1(N924), .B0(n337), .B1(global_cntr[14]), .Y(n39)
         );
  AOI21X1 U48 ( .A0(n626), .A1(\C126/DATA3_15 ), .B0(n41), .Y(\im_a[15]_BAR )
         );
  AO22X1 U49 ( .A0(n356), .A1(N925), .B0(n337), .B1(global_cntr[15]), .Y(n41)
         );
  AOI21X1 U50 ( .A0(n626), .A1(\C126/DATA3_16 ), .B0(n43), .Y(\im_a[16]_BAR )
         );
  AO22X1 U51 ( .A0(n356), .A1(N926), .B0(n337), .B1(global_cntr[16]), .Y(n43)
         );
  AOI21X1 U52 ( .A0(n626), .A1(\C126/DATA3_17 ), .B0(n45), .Y(\im_a[17]_BAR )
         );
  AO22X1 U53 ( .A0(n356), .A1(N927), .B0(n337), .B1(n107), .Y(n45) );
  AOI21X1 U54 ( .A0(n626), .A1(\C126/DATA3_18 ), .B0(n47), .Y(\im_a[18]_BAR )
         );
  AO22X1 U55 ( .A0(n356), .A1(N928), .B0(n337), .B1(global_cntr[18]), .Y(n47)
         );
  AND2X2 U56 ( .A(n252), .B(n377), .Y(n48) );
  OAI2BB2XL U57 ( .B0(n1933), .B1(n1932), .A0N(n1933), .A1N(n49), .Y(n1934) );
  OA22X1 U58 ( .A0(n1789), .A1(n1788), .B0(n1787), .B1(n1786), .Y(n49) );
  NOR2BX1 U59 ( .AN(n1793), .B(n1802), .Y(n1931) );
  AOI2BB1X1 U60 ( .A0N(write_cntr[12]), .A1N(n1206), .B0(n324), .Y(n1219) );
  NAND2X1 U61 ( .A(n902), .B(next_cr_x[5]), .Y(n50) );
  XNOR2X1 U62 ( .A(n50), .B(n903), .Y(n1983) );
  CLKINVX1 U63 ( .A(n511), .Y(n51) );
  CLKINVX1 U64 ( .A(curr_time[1]), .Y(n52) );
  CLKINVX1 U65 ( .A(n528), .Y(n53) );
  AOI221XL U66 ( .A0(n513), .A1(n52), .B0(n520), .B1(curr_time[1]), .C0(n53), 
        .Y(n54) );
  CLKINVX1 U67 ( .A(curr_time[9]), .Y(n55) );
  OAI22XL U68 ( .A0(curr_time[9]), .A1(n512), .B0(n55), .B1(n516), .Y(n56) );
  AO22X1 U69 ( .A0(n514), .A1(n174), .B0(n529), .B1(n56), .Y(n57) );
  AOI211XL U70 ( .A0(n176), .A1(s_1[1]), .B0(n54), .C0(n57), .Y(n58) );
  CLKINVX1 U71 ( .A(n515), .Y(n59) );
  NAND2X1 U72 ( .A(curr_time[17]), .B(n519), .Y(n60) );
  OAI211X1 U73 ( .A0(n59), .A1(curr_time[17]), .B0(n518), .C0(n60), .Y(n61) );
  OAI211X1 U74 ( .A0(n531), .A1(n51), .B0(n58), .C0(n61), .Y(\C1/Z_1 ) );
  CLKINVX1 U75 ( .A(curr_time[7]), .Y(n62) );
  OAI211X1 U76 ( .A0(curr_time[5]), .A1(n62), .B0(n388), .C0(curr_time[6]), 
        .Y(n63) );
  NAND2X1 U77 ( .A(n389), .B(n63), .Y(s_1[3]) );
  NOR2X1 U78 ( .A(n594), .B(n276), .Y(n64) );
  OAI22XL U79 ( .A0(n603), .A1(n2232), .B0(n608), .B1(n539), .Y(n65) );
  AOI211XL U80 ( .A0(n610), .A1(write_addr[17]), .B0(n64), .C0(n65), .Y(n66)
         );
  OAI2BB2XL U81 ( .B0(n618), .B1(n66), .A0N(n48), .A1N(global_cntr[19]), .Y(
        n67) );
  AO22X1 U82 ( .A0(\DP_OP_438J1_134_2124/I5 ), .A1(n67), .B0(si_sel), .B1(N929), .Y(\DP_OP_438J1_134_2124/n64 ) );
  OAI2BB2XL U83 ( .B0(n576), .B1(n266), .A0N(n112), .A1N(n147), .Y(n299) );
  OAI2BB1X1 U84 ( .A0N(n1216), .A1N(n1219), .B0(n1217), .Y(n1281) );
  NAND2BX1 U85 ( .AN(n397), .B(n882), .Y(n456) );
  AOI21X1 U86 ( .A0(next_cr_x[6]), .A1(n710), .B0(n709), .Y(n911) );
  OAI2BB1X1 U87 ( .A0N(n386), .A1N(s_1[3]), .B0(n875), .Y(n395) );
  OAI2BB1X1 U88 ( .A0N(n464), .A1N(n465), .B0(n868), .Y(n475) );
  OAI2BB1X1 U89 ( .A0N(n1248), .A1N(n1250), .B0(n1251), .Y(n1441) );
  CLKINVX1 U90 ( .A(curr_time[23]), .Y(n68) );
  OAI211X1 U91 ( .A0(curr_time[21]), .A1(n68), .B0(n380), .C0(curr_time[22]), 
        .Y(n69) );
  NAND2X1 U92 ( .A(n381), .B(n69), .Y(h_1[3]) );
  NAND2BX1 U93 ( .AN(n169), .B(n1440), .Y(n531) );
  AOI222XL U94 ( .A0(\next_write_addr_w[0] ), .A1(n616), .B0(n632), .B1(n617), 
        .C0(n355), .C1(n615), .Y(n70) );
  OAI22XL U95 ( .A0(n279), .A1(n334), .B0(n618), .B1(n70), .Y(n71) );
  AOI22X1 U96 ( .A0(N910), .A1(si_sel), .B0(\DP_OP_438J1_134_2124/I5 ), .B1(
        n71), .Y(n72) );
  NAND2X1 U97 ( .A(n338), .B(curr_photo_addr[0]), .Y(n73) );
  NOR2X1 U98 ( .A(n72), .B(n73), .Y(\DP_OP_438J1_134_2124/n20 ) );
  AOI2BB2X1 U99 ( .B0(n72), .B1(n73), .A0N(n72), .A1N(n73), .Y(\C126/DATA3_0 )
         );
  AOI2BB2X1 U100 ( .B0(\DP_OP_438J1_134_2124/n64 ), .B1(\C1/Z_19 ), .A0N(
        \DP_OP_438J1_134_2124/n64 ), .A1N(\C1/Z_19 ), .Y(n74) );
  AOI2BB2X1 U101 ( .B0(\DP_OP_438J1_134_2124/n2 ), .B1(n74), .A0N(
        \DP_OP_438J1_134_2124/n2 ), .A1N(n74), .Y(n75) );
  AOI222XL U102 ( .A0(N929), .A1(n356), .B0(n626), .B1(n75), .C0(
        global_cntr[19]), .C1(n337), .Y(\im_a[19]_BAR ) );
  NOR2X1 U103 ( .A(n323), .B(n231), .Y(n76) );
  OA21XL U104 ( .A0(n1951), .A1(n76), .B0(n1942), .Y(n1941) );
  OAI2BB2XL U105 ( .B0(n558), .B1(n266), .A0N(write_addr[13]), .A1N(n147), .Y(
        n294) );
  NOR2X1 U106 ( .A(n708), .B(n219), .Y(n77) );
  XNOR2X1 U107 ( .A(n77), .B(n730), .Y(n743) );
  NAND2X1 U108 ( .A(n2004), .B(n2156), .Y(n78) );
  XNOR2X1 U109 ( .A(n78), .B(n786), .Y(n799) );
  OAI2BB1X1 U110 ( .A0N(n1229), .A1N(n1232), .B0(n1230), .Y(n1280) );
  XNOR2X1 U111 ( .A(n809), .B(n808), .Y(n164) );
  NOR2X1 U112 ( .A(n180), .B(next_cr_x[5]), .Y(n79) );
  OAI21XL U113 ( .A0(n79), .A1(n1993), .B0(n1976), .Y(n80) );
  XNOR2X1 U114 ( .A(n1977), .B(n80), .Y(n1992) );
  CLKINVX1 U115 ( .A(curr_time[12]), .Y(n81) );
  NAND2X1 U116 ( .A(n467), .B(n475), .Y(n82) );
  OAI211X1 U117 ( .A0(n868), .A1(n81), .B0(n870), .C0(n82), .Y(n474) );
  CLKINVX1 U118 ( .A(curr_time[2]), .Y(n83) );
  AO21X1 U119 ( .A0(n83), .A1(s_1[1]), .B0(n881), .Y(n459) );
  AO21X1 U120 ( .A0(\DP_OP_166J1_126_2191/n24 ), .A1(n179), .B0(
        \DP_OP_166J1_126_2191/I2 ), .Y(n84) );
  AND2X1 U121 ( .A(\DP_OP_166J1_126_2191/n4 ), .B(n84), .Y(
        \DP_OP_166J1_126_2191/n3 ) );
  AOI2BB2X1 U122 ( .B0(\DP_OP_166J1_126_2191/n4 ), .B1(n84), .A0N(
        \DP_OP_166J1_126_2191/n4 ), .A1N(n84), .Y(N689) );
  NOR3X1 U123 ( .A(n279), .B(global_cntr[1]), .C(n1283), .Y(N1571) );
  NAND3BX1 U124 ( .AN(n1933), .B(n26), .C(en_so), .Y(n85) );
  CLKINVX1 U125 ( .A(n85), .Y(n632) );
  OAI2BB2XL U126 ( .B0(n2229), .B1(n266), .A0N(write_addr[11]), .A1N(n147), 
        .Y(n296) );
  OAI2BB1X1 U127 ( .A0N(n754), .A1N(n751), .B0(n756), .Y(n2140) );
  OAI2BB1X1 U128 ( .A0N(n1244), .A1N(n1246), .B0(n1245), .Y(n1279) );
  OAI2BB1X1 U129 ( .A0N(n378), .A1N(h_1[3]), .B0(n860), .Y(n434) );
  NAND2X1 U130 ( .A(n1979), .B(n2107), .Y(n86) );
  XNOR2X1 U131 ( .A(n86), .B(n1980), .Y(n1990) );
  OAI2BB1X1 U132 ( .A0N(n1639), .A1N(n1644), .B0(n1636), .Y(n1637) );
  CLKINVX1 U133 ( .A(curr_time[4]), .Y(n87) );
  NAND2X1 U134 ( .A(n389), .B(n395), .Y(n88) );
  OAI211X1 U135 ( .A0(n875), .A1(n87), .B0(n876), .C0(n88), .Y(n394) );
  CLKINVX1 U136 ( .A(curr_time[14]), .Y(n89) );
  OA21XL U137 ( .A0(n466), .A1(n89), .B0(n467), .Y(n476) );
  OAI2BB1X1 U138 ( .A0N(n709), .A1N(n710), .B0(n728), .Y(n718) );
  AOI2BB1X1 U139 ( .A0N(n816), .A1N(n814), .B0(n810), .Y(n2167) );
  XNOR2X1 U140 ( .A(n921), .B(n920), .Y(n923) );
  AOI2BB2X1 U141 ( .B0(write_addr[19]), .B1(fb_addr[19]), .A0N(write_addr[19]), 
        .A1N(fb_addr[19]), .Y(n90) );
  AOI2BB2X1 U142 ( .B0(\DP_OP_438J1_134_2124/n22 ), .B1(n90), .A0N(
        \DP_OP_438J1_134_2124/n22 ), .A1N(n90), .Y(N929) );
  AO21X1 U143 ( .A0(\DP_OP_166J1_126_2191/n25 ), .A1(n179), .B0(
        \DP_OP_166J1_126_2191/I2 ), .Y(n91) );
  AND2X1 U144 ( .A(\DP_OP_166J1_126_2191/n3 ), .B(n91), .Y(
        \DP_OP_166J1_126_2191/n2 ) );
  AOI2BB2X1 U145 ( .B0(\DP_OP_166J1_126_2191/n3 ), .B1(n91), .A0N(
        \DP_OP_166J1_126_2191/n3 ), .A1N(n91), .Y(N690) );
  AND3X1 U146 ( .A(global_cntr[7]), .B(global_cntr[6]), .C(n652), .Y(n365) );
  NAND3X1 U147 ( .A(n1282), .B(n657), .C(n226), .Y(n92) );
  NOR2X1 U148 ( .A(N1593), .B(n92), .Y(en_fb_addr) );
  OAI2BB2XL U149 ( .B0(n593), .B1(n266), .A0N(write_addr[4]), .A1N(n147), .Y(
        n303) );
  NAND2BX1 U150 ( .AN(n2134), .B(n2136), .Y(n2141) );
  CLKINVX1 U151 ( .A(curr_time[20]), .Y(n93) );
  NAND2X1 U152 ( .A(n381), .B(n434), .Y(n94) );
  OAI211X1 U153 ( .A0(n860), .A1(n93), .B0(n863), .C0(n94), .Y(n433) );
  AO22X1 U154 ( .A0(n95), .A1(n1245), .B0(n1246), .B1(n1244), .Y(n1251) );
  CLKINVX1 U155 ( .A(n1246), .Y(n95) );
  OAI2BB1X1 U156 ( .A0N(n479), .A1N(n484), .B0(n485), .Y(n511) );
  CLKINVX1 U157 ( .A(n658), .Y(n96) );
  AOI2BB2X1 U158 ( .B0(n96), .B1(n883), .A0N(n96), .A1N(s_1[1]), .Y(n884) );
  NAND2X1 U159 ( .A(n1991), .B(n2095), .Y(n97) );
  XNOR2X1 U160 ( .A(n97), .B(n1992), .Y(n2012) );
  CLKINVX1 U161 ( .A(n2170), .Y(n98) );
  CLKINVX1 U162 ( .A(n2171), .Y(n99) );
  OAI32X1 U163 ( .A0(n2171), .A1(n2169), .A2(n98), .B0(n2170), .B1(n99), .Y(
        n2180) );
  CLKINVX1 U164 ( .A(n919), .Y(n100) );
  OAI211X1 U165 ( .A0(n921), .A1(n920), .B0(n322), .C0(n100), .Y(n101) );
  NAND2X1 U166 ( .A(n922), .B(n101), .Y(n535) );
  AOI2BB2X1 U167 ( .B0(n170), .B1(next_cr_x[5]), .A0N(n170), .A1N(next_cr_x[5]), .Y(n102) );
  AOI2BB2X1 U168 ( .B0(n102), .B1(next_cr_x[6]), .A0N(n102), .A1N(next_cr_x[6]), .Y(\DP_OP_436J1_125_1438/n26 ) );
  NAND3BX1 U169 ( .AN(n704), .B(write_cntr[12]), .C(write_cntr[13]), .Y(n702)
         );
  OAI2BB1X1 U170 ( .A0N(n1658), .A1N(n1663), .B0(n1655), .Y(n1656) );
  AO21X1 U171 ( .A0(\DP_OP_166J1_126_2191/n26 ), .A1(n179), .B0(
        \DP_OP_166J1_126_2191/I2 ), .Y(n103) );
  AND2X1 U172 ( .A(\DP_OP_166J1_126_2191/n2 ), .B(n103), .Y(
        \DP_OP_166J1_126_2191/n1 ) );
  AOI2BB2X1 U173 ( .B0(\DP_OP_166J1_126_2191/n2 ), .B1(n103), .A0N(
        \DP_OP_166J1_126_2191/n2 ), .A1N(n103), .Y(N691) );
  NAND2X1 U174 ( .A(n2214), .B(n421), .Y(n104) );
  OAI211X1 U175 ( .A0(n2214), .A1(n421), .B0(n660), .C0(n104), .Y(n539) );
  OAI2BB1X1 U176 ( .A0N(n1493), .A1N(n1494), .B0(n1495), .Y(n105) );
  NAND2X1 U177 ( .A(n105), .B(n1498), .Y(n1496) );
  AOI21X1 U178 ( .A0(n331), .A1(n2222), .B0(n2221), .Y(next_photo[0]) );
  AOI2BB1X1 U179 ( .A0N(n648), .A1N(global_cntr[10]), .B0(n366), .Y(n647) );
  AO21X1 U180 ( .A0(n106), .A1(n657), .B0(n924), .Y(next_glb_cntr[2]) );
  CLKINVX1 U181 ( .A(global_cntr[2]), .Y(n106) );
  OAI2BB2XL U182 ( .B0(n2233), .B1(n147), .A0N(write_addr[3]), .A1N(n266), .Y(
        n304) );
  CLKINVX1 U183 ( .A(n2049), .Y(n171) );
  BUFX4 U184 ( .A(n359), .Y(n358) );
  CLKBUFX3 U185 ( .A(n114), .Y(n359) );
  NOR2X2 U186 ( .A(n227), .B(n257), .Y(n1911) );
  CLKINVX1 U187 ( .A(n320), .Y(n107) );
  INVXL U188 ( .A(n322), .Y(n108) );
  CLKBUFX2 U189 ( .A(write_addr[9]), .Y(n109) );
  CLKINVX1 U190 ( .A(n327), .Y(n110) );
  INVXL U191 ( .A(n256), .Y(n111) );
  CLKINVX1 U192 ( .A(n278), .Y(n112) );
  NOR2X1 U193 ( .A(N76), .B(N1182), .Y(n1427) );
  INVXL U194 ( .A(write_cntr[10]), .Y(n113) );
  NOR2X2 U195 ( .A(work_cntr[19]), .B(n236), .Y(n1798) );
  AOI2BB2X2 U196 ( .B0(work_cntr[13]), .B1(n1320), .A0N(work_cntr[13]), .A1N(
        n1320), .Y(n1318) );
  NAND2X2 U197 ( .A(N76), .B(N1182), .Y(n1189) );
  OAI21X4 U198 ( .A0(N76), .A1(N1182), .B0(n1189), .Y(n1778) );
  OAI21X2 U199 ( .A0(n1108), .A1(n267), .B0(n1107), .Y(n1129) );
  AOI2BB2X2 U200 ( .B0(n947), .B1(n264), .A0N(n947), .A1N(n264), .Y(n951) );
  INVX6 U201 ( .A(reset), .Y(n114) );
  CLKINVX1 U234 ( .A(im_wen_n), .Y(n420) );
  AND3X2 U235 ( .A(n169), .B(n525), .C(n524), .Y(\DP_OP_166J1_126_2191/I2 ) );
  NOR2X2 U236 ( .A(n454), .B(n525), .Y(n528) );
  AND2X2 U237 ( .A(n2135), .B(n2134), .Y(n237) );
  BUFX2 U238 ( .A(n2023), .Y(n177) );
  OR2XL U239 ( .A(N76), .B(n149), .Y(next_work_cntr[0]) );
  OAI21X1 U240 ( .A0(n267), .A1(n979), .B0(n977), .Y(n985) );
  NAND2X1 U241 ( .A(n656), .B(n1614), .Y(n2218) );
  OAI22X1 U242 ( .A0(n1620), .A1(n1619), .B0(n1618), .B1(work_cntr[19]), .Y(
        n1629) );
  CLKINVX1 U243 ( .A(n1625), .Y(n148) );
  NOR2X1 U244 ( .A(global_cntr[6]), .B(global_cntr[12]), .Y(n930) );
  OA21XL U245 ( .A0(n856), .A1(n855), .B0(n854), .Y(\next_cr_y[0] ) );
  OAI221X1 U246 ( .A0(n1572), .A1(n1574), .B0(n1571), .B1(n1570), .C0(n1569), 
        .Y(n1578) );
  NOR2X2 U247 ( .A(n818), .B(n823), .Y(n2172) );
  AOI31X1 U248 ( .A0(n813), .A1(n812), .A2(n2170), .B0(n811), .Y(n830) );
  OA21XL U249 ( .A0(n1762), .A1(n1761), .B0(n1760), .Y(n1770) );
  OAI31X1 U250 ( .A0(n817), .A1(n2167), .A2(n816), .B0(n815), .Y(n823) );
  OAI31X1 U251 ( .A0(n1425), .A1(n1424), .A2(n1423), .B0(n1422), .Y(n1433) );
  AOI211X1 U252 ( .A0(n257), .A1(n1419), .B0(n1423), .C0(n1408), .Y(n1411) );
  OAI31X1 U253 ( .A0(n1515), .A1(n1514), .A2(n1513), .B0(n1512), .Y(n1520) );
  OAI21XL U254 ( .A0(n1731), .A1(n1733), .B0(n1730), .Y(n1743) );
  OA21XL U255 ( .A0(n1723), .A1(n1722), .B0(n1721), .Y(n1729) );
  OA22XL U256 ( .A0(n1997), .A1(n2088), .B0(n2004), .B1(n2095), .Y(n2025) );
  OAI31X1 U257 ( .A0(n1498), .A1(n1497), .A2(n1506), .B0(n1496), .Y(n1500) );
  OAI211X1 U258 ( .A0(n1542), .A1(n1394), .B0(n1391), .C0(n1395), .Y(n1392) );
  OAI31X1 U259 ( .A0(n1708), .A1(n1707), .A2(n1706), .B0(n1705), .Y(n1715) );
  AOI221X1 U260 ( .A0(n1504), .A1(n1502), .B0(n1501), .B1(n1502), .C0(n1503), 
        .Y(n1506) );
  AND3X2 U261 ( .A(n533), .B(n532), .C(n531), .Y(\DP_OP_166J1_126_2191/I3 ) );
  OA21XL U262 ( .A0(n1703), .A1(n1702), .B0(n1701), .Y(n1709) );
  OA21XL U263 ( .A0(n1026), .A1(n1030), .B0(n1025), .Y(n1032) );
  OR2XL U264 ( .A(n490), .B(n525), .Y(n527) );
  AND3X2 U265 ( .A(n490), .B(n155), .C(n453), .Y(n526) );
  OAI31X1 U266 ( .A0(n744), .A1(n743), .A2(n742), .B0(n741), .Y(n754) );
  OR2XL U267 ( .A(n1441), .B(n524), .Y(n530) );
  OAI211X1 U268 ( .A0(n1471), .A1(n173), .B0(n1472), .C0(n1469), .Y(n1478) );
  OA21XL U269 ( .A0(n1356), .A1(n1355), .B0(n1357), .Y(n1378) );
  OA21XL U270 ( .A0(n1683), .A1(n1682), .B0(n1681), .Y(n1689) );
  OAI31X1 U271 ( .A0(n1351), .A1(n1350), .A2(n1349), .B0(n1348), .Y(n1356) );
  AOI222X1 U272 ( .A0(n712), .A1(n2087), .B0(n712), .B1(n711), .C0(n710), .C1(
        next_cr_x[6]), .Y(n901) );
  AOI2BB2X1 U273 ( .B0(n1463), .B1(n1462), .A0N(n1463), .A1N(n1462), .Y(n1467)
         );
  OAI31X1 U274 ( .A0(n994), .A1(work_cntr[9]), .A2(n993), .B0(n992), .Y(n999)
         );
  OA21XL U275 ( .A0(n1663), .A1(n1662), .B0(n1661), .Y(n1669) );
  OR2X2 U276 ( .A(n217), .B(n218), .Y(n216) );
  OA21XL U277 ( .A0(n1143), .A1(n1142), .B0(n1141), .Y(n1146) );
  OAI211X1 U278 ( .A0(n2210), .A1(n2209), .B0(n660), .C0(n2212), .Y(n2232) );
  OAI211X1 U279 ( .A0(n2207), .A1(n2206), .B0(n660), .C0(n2208), .Y(n2231) );
  INVX6 U280 ( .A(n220), .Y(n149) );
  OAI211X1 U281 ( .A0(n334), .A1(n692), .B0(n685), .C0(n684), .Y(n689) );
  CLKINVX1 U282 ( .A(n171), .Y(n150) );
  NOR2BX1 U283 ( .AN(n686), .B(n2241), .Y(n376) );
  OAI211X1 U284 ( .A0(n1290), .A1(n1293), .B0(n1292), .C0(n1297), .Y(n1304) );
  AOI211X1 U285 ( .A0(n247), .A1(n373), .B0(n664), .C0(n375), .Y(n639) );
  OR2X1 U286 ( .A(n212), .B(n213), .Y(n211) );
  OR2XL U287 ( .A(n222), .B(n1627), .Y(n1625) );
  OAI211X1 U288 ( .A0(n923), .A1(n322), .B0(n538), .C0(n534), .Y(n536) );
  OR2X1 U289 ( .A(n205), .B(n206), .Y(n204) );
  OA21XL U290 ( .A0(n1886), .A1(n229), .B0(n1885), .Y(n1902) );
  NAND2X1 U291 ( .A(n26), .B(n1936), .Y(n1435) );
  INVX6 U292 ( .A(n2241), .Y(si_sel) );
  NAND2BX2 U293 ( .AN(n932), .B(n26), .Y(N1593) );
  NAND2X1 U294 ( .A(curr_time[23]), .B(n859), .Y(n381) );
  NOR2X1 U295 ( .A(curr_time[21]), .B(curr_time[22]), .Y(n859) );
  NAND2X1 U296 ( .A(n790), .B(n789), .Y(n793) );
  NAND2BX1 U297 ( .AN(n954), .B(n953), .Y(n958) );
  CLKINVX1 U298 ( .A(n1743), .Y(n152) );
  OA21X1 U299 ( .A0(n265), .A1(n998), .B0(n997), .Y(n1004) );
  NAND2BX1 U300 ( .AN(n1913), .B(n1910), .Y(n1920) );
  NAND2X1 U301 ( .A(n732), .B(n731), .Y(n735) );
  CLKINVX1 U302 ( .A(n729), .Y(n732) );
  NAND2X1 U303 ( .A(n1447), .B(n730), .Y(n731) );
  NOR2X2 U304 ( .A(n149), .B(n1711), .Y(next_work_cntr[8]) );
  NOR2X1 U305 ( .A(n657), .B(n226), .Y(n924) );
  AOI211X1 U306 ( .A0(n1200), .A1(n1199), .B0(n2225), .C0(n1198), .Y(n2224) );
  CLKINVX1 U307 ( .A(n2236), .Y(n2225) );
  NOR2X1 U308 ( .A(n2087), .B(n2088), .Y(n2111) );
  INVXL U309 ( .A(next_work_cntr[0]), .Y(n153) );
  MXI2X2 U310 ( .A(n332), .B(n333), .S0(next_cr_x[5]), .Y(
        \DP_OP_436J1_125_1438/n25 ) );
  NAND3X1 U311 ( .A(n1167), .B(n1166), .C(n1168), .Y(n1180) );
  NOR2X1 U312 ( .A(n2088), .B(n2004), .Y(n2003) );
  INVX3 U313 ( .A(n2095), .Y(n2088) );
  NOR2X1 U314 ( .A(n273), .B(n2115), .Y(n2126) );
  OAI21X1 U315 ( .A0(n1868), .A1(n1867), .B0(n1866), .Y(n1871) );
  OAI21X1 U316 ( .A0(n1803), .A1(n260), .B0(n1802), .Y(n1805) );
  OAI21X1 U317 ( .A0(n2200), .A1(n2204), .B0(n2199), .Y(n2201) );
  NAND4X1 U318 ( .A(n109), .B(n110), .C(write_addr[12]), .D(n2198), .Y(n2204)
         );
  INVXL U319 ( .A(n633), .Y(n154) );
  CLKINVX1 U320 ( .A(n154), .Y(n155) );
  OAI21X1 U321 ( .A0(n1777), .A1(n1776), .B0(n1778), .Y(n1780) );
  OAI21X1 U322 ( .A0(n229), .A1(n1031), .B0(n1030), .Y(n1034) );
  OAI21X1 U323 ( .A0(n1756), .A1(n1764), .B0(n1761), .Y(n1757) );
  OAI21X1 U324 ( .A0(n1644), .A1(n1643), .B0(n1642), .Y(n1650) );
  INVXL U325 ( .A(n1669), .Y(n156) );
  INVXL U326 ( .A(n1689), .Y(n157) );
  INVXL U327 ( .A(n1709), .Y(n158) );
  INVXL U328 ( .A(n1729), .Y(n159) );
  OAI21X1 U329 ( .A0(n1010), .A1(n1014), .B0(n1009), .Y(n1016) );
  INVXL U330 ( .A(n1032), .Y(n160) );
  INVXL U331 ( .A(n1770), .Y(n161) );
  AOI21X1 U332 ( .A0(n1496), .A1(n1491), .B0(n1490), .Y(n1492) );
  OAI21X1 U333 ( .A0(n1048), .A1(n1049), .B0(n1047), .Y(n1051) );
  AOI31X1 U334 ( .A0(n1370), .A1(n1362), .A2(n1361), .B0(n1360), .Y(n1364) );
  OAI21X1 U335 ( .A0(n1881), .A1(n1880), .B0(n1879), .Y(n1884) );
  INVXL U336 ( .A(n1146), .Y(n162) );
  CLKINVX1 U337 ( .A(n2025), .Y(n163) );
  AOI32X1 U338 ( .A0(n220), .A1(n702), .A2(write_cntr[13]), .B0(n703), .B1(
        n702), .Y(n729) );
  OAI21X1 U339 ( .A0(n1768), .A1(n1772), .B0(n1767), .Y(n1775) );
  OAI21X1 U340 ( .A0(n1296), .A1(n1295), .B0(n1294), .Y(n1300) );
  AOI32X1 U341 ( .A0(n1626), .A1(n940), .A2(n260), .B0(n941), .B1(n940), .Y(
        n942) );
  INVXL U342 ( .A(n1211), .Y(n165) );
  CLKINVX1 U343 ( .A(n165), .Y(n166) );
  AOI2BB2X2 U344 ( .B0(n1223), .B1(n1222), .A0N(n1223), .A1N(n1222), .Y(n1241)
         );
  OAI22X1 U345 ( .A0(n1316), .A1(n1315), .B0(n1314), .B1(n1313), .Y(n1317) );
  INVXL U346 ( .A(n1755), .Y(n167) );
  INVXL U347 ( .A(n167), .Y(n168) );
  AOI211X1 U348 ( .A0(n660), .A1(n1936), .B0(n1939), .C0(n659), .Y(n2243) );
  AOI31X1 U349 ( .A0(work_cntr[4]), .A1(n220), .A2(n1457), .B0(
        next_work_cntr[5]), .Y(n1545) );
  NOR3X1 U350 ( .A(n230), .B(n248), .C(n221), .Y(n1203) );
  OAI21X1 U351 ( .A0(n906), .A1(n1976), .B0(n905), .Y(n907) );
  NAND2X1 U352 ( .A(n180), .B(next_cr_x[5]), .Y(n1976) );
  OAI21X1 U353 ( .A0(n1237), .A1(n1257), .B0(n1236), .Y(n1238) );
  AOI211X1 U354 ( .A0(n1563), .A1(n1561), .B0(n1569), .C0(n1560), .Y(n1575) );
  OAI31X1 U355 ( .A0(n2027), .A1(n2030), .A2(n2032), .B0(n2035), .Y(n2034) );
  NOR2X2 U356 ( .A(n935), .B(n259), .Y(n1792) );
  NOR2X1 U357 ( .A(n365), .B(n364), .Y(n651) );
  OAI31X1 U358 ( .A0(n754), .A1(n2138), .A2(n753), .B0(n752), .Y(n760) );
  OAI2BB2X1 U359 ( .B0(n1161), .B1(n1160), .A0N(n1161), .A1N(n1159), .Y(n1170)
         );
  NOR2X1 U360 ( .A(n149), .B(N1184), .Y(n1585) );
  OAI21X1 U361 ( .A0(n652), .A1(n246), .B0(n363), .Y(next_glb_cntr[6]) );
  OAI21X1 U362 ( .A0(n2217), .A1(n2216), .B0(n2215), .Y(n2222) );
  NOR2X1 U363 ( .A(n1427), .B(n257), .Y(n2237) );
  NOR2X1 U364 ( .A(n851), .B(n850), .Y(n2039) );
  CLKINVX1 U365 ( .A(n2124), .Y(n850) );
  OAI31X1 U366 ( .A0(n1263), .A1(n1262), .A2(n1271), .B0(n1276), .Y(n1438) );
  NOR4X1 U367 ( .A(n1268), .B(n1264), .C(n1267), .D(n285), .Y(n1263) );
  NAND2X1 U368 ( .A(n1356), .B(n1355), .Y(n1368) );
  OAI21X1 U369 ( .A0(n1863), .A1(n265), .B0(n1847), .Y(n1355) );
  NOR2X1 U370 ( .A(n261), .B(n885), .Y(n888) );
  OAI211X1 U371 ( .A0(n2150), .A1(n2152), .B0(n2149), .C0(n2148), .Y(n2155) );
  OAI21X1 U372 ( .A0(n2144), .A1(n2143), .B0(n2142), .Y(n2150) );
  OAI31X1 U373 ( .A0(n1021), .A1(work_cntr[6]), .A2(n1020), .B0(n1019), .Y(
        n1028) );
  OAI21X1 U374 ( .A0(n261), .A1(n1015), .B0(n1014), .Y(n1020) );
  OAI2BB2X1 U375 ( .B0(work_cntr[6]), .B1(n1791), .A0N(work_cntr[6]), .A1N(
        n1791), .Y(n1384) );
  OAI21X1 U376 ( .A0(n1060), .A1(n1059), .B0(n1058), .Y(n1063) );
  OAI21X1 U377 ( .A0(n1451), .A1(n1188), .B0(n1196), .Y(n1197) );
  OAI21X1 U378 ( .A0(n747), .A1(n746), .B0(n745), .Y(n756) );
  OAI22X1 U379 ( .A0(n1243), .A1(n1242), .B0(n1245), .B1(n1244), .Y(n1248) );
  NAND2X1 U380 ( .A(curr_time[15]), .B(n867), .Y(n467) );
  NAND2X1 U381 ( .A(curr_time[7]), .B(n874), .Y(n389) );
  NOR2X1 U382 ( .A(curr_time[17]), .B(n515), .Y(n497) );
  AOI22X1 U383 ( .A0(\DP_OP_436J1_125_1438/n26 ), .A1(n659), .B0(n2104), .B1(
        n2103), .Y(n576) );
  NOR2X2 U384 ( .A(n695), .B(n696), .Y(n2104) );
  CLKINVX1 U385 ( .A(n219), .Y(n2134) );
  CLKINVX1 U386 ( .A(n2185), .Y(n2179) );
  OAI21X1 U387 ( .A0(work_cntr[18]), .A1(n148), .B0(n1623), .Y(n1621) );
  AOI22X1 U388 ( .A0(n1623), .A1(work_cntr[19]), .B0(n1798), .B1(n148), .Y(
        n1456) );
  CLKINVX1 U389 ( .A(curr_time[10]), .Y(n482) );
  NAND2X1 U390 ( .A(work_cntr[18]), .B(n148), .Y(n1623) );
  OAI21X1 U391 ( .A0(n511), .A1(n482), .B0(n483), .Y(n504) );
  NAND2X1 U392 ( .A(n511), .B(n482), .Y(n483) );
  NAND2X1 U393 ( .A(n1463), .B(n1462), .Y(n1596) );
  CLKINVX1 U394 ( .A(next_work_cntr[18]), .Y(n1463) );
  NOR2X1 U395 ( .A(n1912), .B(n1911), .Y(n1916) );
  NOR2X1 U396 ( .A(n286), .B(n1950), .Y(n1954) );
  AND2X2 U397 ( .A(global_cntr[1]), .B(global_cntr[0]), .Y(n657) );
  OAI31X1 U398 ( .A0(global_cntr[0]), .A1(n249), .A2(n226), .B0(n1614), .Y(
        n692) );
  NAND2X1 U399 ( .A(n1771), .B(n1773), .Y(n1784) );
  NAND2X1 U400 ( .A(n1637), .B(n1638), .Y(n1649) );
  NAND2X1 U401 ( .A(n515), .B(n438), .Y(n519) );
  NAND2X1 U402 ( .A(n1656), .B(n1657), .Y(n1668) );
  NAND2X1 U403 ( .A(n1013), .B(n1015), .Y(n1021) );
  NAND2X1 U404 ( .A(n1696), .B(n1697), .Y(n1708) );
  NAND2X1 U405 ( .A(n1676), .B(n1677), .Y(n1688) );
  CLKINVX1 U406 ( .A(n852), .Y(n2042) );
  NAND2X1 U407 ( .A(n1716), .B(n1717), .Y(n1728) );
  CLKINVX1 U408 ( .A(n1177), .Y(n1182) );
  AND2X2 U409 ( .A(n470), .B(n469), .Y(n487) );
  NAND2X1 U410 ( .A(n1413), .B(n1284), .Y(n1426) );
  CLKINVX1 U411 ( .A(n177), .Y(n1445) );
  AOI32X1 U412 ( .A0(n1815), .A1(n1814), .A2(n1813), .B0(n1812), .B1(n1814), 
        .Y(n1818) );
  NAND2X1 U413 ( .A(n1804), .B(n1812), .Y(n1814) );
  NOR2BX1 U414 ( .AN(n1368), .B(n1360), .Y(n1357) );
  CLKINVX1 U415 ( .A(n1254), .Y(n1267) );
  NOR2X1 U416 ( .A(n1257), .B(n1255), .Y(n1254) );
  NAND2X1 U417 ( .A(n1083), .B(n1093), .Y(n1092) );
  NOR2X1 U418 ( .A(n2081), .B(n239), .Y(n1963) );
  XNOR2X1 U419 ( .A(n2081), .B(write_addr[5]), .Y(n630) );
  NAND2X1 U420 ( .A(n2080), .B(write_addr[4]), .Y(n2081) );
  CLKINVX1 U421 ( .A(n748), .Y(n759) );
  OAI31X1 U422 ( .A0(n759), .A1(n758), .A2(n2138), .B0(n757), .Y(n771) );
  CLKINVX1 U423 ( .A(n532), .Y(n518) );
  NOR2X1 U424 ( .A(n759), .B(n758), .Y(n751) );
  NAND2X1 U425 ( .A(n1495), .B(n1494), .Y(n1503) );
  NOR2X1 U426 ( .A(n1490), .B(n1497), .Y(n1495) );
  CLKINVX1 U427 ( .A(next_work_cntr[13]), .Y(n1487) );
  NOR2X1 U428 ( .A(n149), .B(n1658), .Y(next_work_cntr[13]) );
  NOR2X1 U429 ( .A(n2050), .B(n2052), .Y(n2053) );
  NOR2X1 U430 ( .A(n2212), .B(n321), .Y(n421) );
  AOI211X1 U431 ( .A0(n2212), .A1(n2213), .B0(n2211), .C0(n421), .Y(n540) );
  NAND2X1 U432 ( .A(n2210), .B(n2209), .Y(n2212) );
  NAND2X1 U433 ( .A(n1249), .B(n1441), .Y(n1260) );
  NOR3X2 U434 ( .A(n2203), .B(n274), .C(n2199), .Y(n1957) );
  NAND2BX1 U435 ( .AN(n1045), .B(n1050), .Y(n1057) );
  NAND2X1 U436 ( .A(n1235), .B(n1236), .Y(n1259) );
  NAND2X1 U437 ( .A(global_cntr[13]), .B(n368), .Y(n369) );
  AOI211X1 U438 ( .A0(n243), .A1(n369), .B0(n370), .C0(n375), .Y(n643) );
  OA21XL U439 ( .A0(global_cntr[11]), .A1(n366), .B0(n367), .Y(n646) );
  AND2X2 U440 ( .A(n648), .B(global_cntr[10]), .Y(n366) );
  INVXL U441 ( .A(n526), .Y(n169) );
  NAND2X1 U442 ( .A(n25), .B(n24), .Y(n932) );
  NAND2X1 U443 ( .A(n234), .B(n25), .Y(n687) );
  NOR2X1 U444 ( .A(n234), .B(n25), .Y(n694) );
  NAND2X1 U445 ( .A(write_addr[11]), .B(n2174), .Y(n2187) );
  NAND2BX1 U446 ( .AN(n2211), .B(n418), .Y(n550) );
  NAND2X1 U447 ( .A(n1337), .B(n1336), .Y(n1342) );
  CLKINVX1 U448 ( .A(n1523), .Y(n1518) );
  NAND2X1 U449 ( .A(n1517), .B(n1516), .Y(n1523) );
  AND2X2 U450 ( .A(n2179), .B(n2178), .Y(n232) );
  ADDFX2 U451 ( .A(n2118), .B(n2133), .CI(n2132), .CO(n2178), .S(n2131) );
  NAND2X1 U452 ( .A(n1224), .B(n1280), .Y(n1227) );
  NAND2BX1 U453 ( .AN(n2211), .B(n419), .Y(n554) );
  NOR2BX1 U454 ( .AN(n2199), .B(n2200), .Y(n2191) );
  AOI2BB2X2 U455 ( .B0(next_work_cntr[14]), .B1(n1475), .A0N(
        next_work_cntr[14]), .A1N(n1475), .Y(n1485) );
  NAND2X1 U456 ( .A(n1486), .B(n1487), .Y(n1475) );
  NAND2X1 U457 ( .A(n1968), .B(write_addr[8]), .Y(n2115) );
  CLKINVX1 U458 ( .A(n1964), .Y(n1968) );
  AOI2BB2X2 U459 ( .B0(n1466), .B1(next_work_cntr[15]), .A0N(n1466), .A1N(
        next_work_cntr[15]), .Y(n1480) );
  NOR2X1 U460 ( .A(n1475), .B(next_work_cntr[14]), .Y(n1466) );
  OAI22X1 U461 ( .A0(n178), .A1(n1901), .B0(n1900), .B1(n1899), .Y(n1914) );
  NOR2BX1 U462 ( .AN(n1898), .B(n1897), .Y(n1900) );
  OAI21X1 U463 ( .A0(n1969), .A1(n276), .B0(n1968), .Y(n1972) );
  XNOR2X1 U464 ( .A(write_addr[19]), .B(n1969), .Y(n2214) );
  NAND2X1 U465 ( .A(n1962), .B(write_addr[18]), .Y(n1969) );
  NAND2X1 U466 ( .A(n487), .B(n482), .Y(n484) );
  OAI22X1 U467 ( .A0(n1112), .A1(n1104), .B0(n1103), .B1(n1102), .Y(n1113) );
  NOR2BX1 U468 ( .AN(n1098), .B(n1089), .Y(n1103) );
  ADDFX2 U469 ( .A(n2107), .B(n2106), .CI(n2105), .CO(n2109), .S(n2098) );
  NOR2X1 U470 ( .A(n2082), .B(n2083), .Y(n2106) );
  NOR2X1 U471 ( .A(n2092), .B(n2078), .Y(n2094) );
  NAND2BX1 U472 ( .AN(n960), .B(n962), .Y(n969) );
  OAI31X1 U473 ( .A0(n969), .A1(work_cntr[12]), .A2(n968), .B0(n967), .Y(n976)
         );
  NAND2BX1 U474 ( .AN(n983), .B(n984), .Y(n994) );
  OAI31X1 U475 ( .A0(n1402), .A1(n1401), .A2(n1400), .B0(n1399), .Y(n1403) );
  NOR2X1 U476 ( .A(n1405), .B(n1404), .Y(n1400) );
  NAND3X1 U477 ( .A(n1440), .B(n453), .C(n1441), .Y(n525) );
  NOR2X1 U478 ( .A(n639), .B(n638), .Y(n678) );
  NOR2X1 U479 ( .A(n270), .B(n821), .Y(n807) );
  NAND2X1 U480 ( .A(cr_read_cntr[8]), .B(n287), .Y(n914) );
  NAND2X1 U481 ( .A(n827), .B(n820), .Y(n834) );
  NOR2X1 U482 ( .A(n2088), .B(n2072), .Y(n2085) );
  NAND2BX1 U483 ( .AN(n836), .B(n1443), .Y(n840) );
  NAND2X1 U484 ( .A(n700), .B(n699), .Y(n1940) );
  NOR2X2 U485 ( .A(n2069), .B(n2060), .Y(n2059) );
  NOR2X1 U486 ( .A(n2058), .B(n2071), .Y(n2069) );
  AOI2BB2X2 U487 ( .B0(work_cntr[7]), .B1(n1285), .A0N(work_cntr[7]), .A1N(
        n1285), .Y(n1375) );
  NAND2X1 U488 ( .A(n1791), .B(n263), .Y(n1285) );
  NAND2BX1 U489 ( .AN(n972), .B(n971), .Y(n975) );
  NOR2X1 U490 ( .A(n964), .B(n963), .Y(n972) );
  NAND2X1 U491 ( .A(write_cntr[14]), .B(n1204), .Y(n1217) );
  NAND2X1 U492 ( .A(global_cntr[11]), .B(n366), .Y(n367) );
  NAND2BX1 U493 ( .AN(n1635), .B(n1634), .Y(n1641) );
  NOR2X1 U494 ( .A(n1624), .B(n1630), .Y(n1635) );
  NOR2X1 U495 ( .A(n837), .B(n716), .Y(n707) );
  AOI21X1 U496 ( .A0(write_cntr[4]), .A1(n1440), .B0(n1264), .Y(n1269) );
  NAND2BX1 U497 ( .AN(n1323), .B(n1319), .Y(n1324) );
  NOR2X1 U498 ( .A(cr_read_cntr[5]), .B(n917), .Y(n919) );
  NOR2X1 U499 ( .A(n1485), .B(n1483), .Y(n1497) );
  OAI2BB2X1 U500 ( .B0(n1482), .B1(n1481), .A0N(n1480), .A1N(n1479), .Y(n1483)
         );
  OAI2BB2X1 U501 ( .B0(next_work_cntr[8]), .B1(n1536), .A0N(next_work_cntr[8]), 
        .A1N(n1536), .Y(n1548) );
  NOR2X1 U502 ( .A(n1305), .B(n1314), .Y(n1311) );
  NOR2BX1 U503 ( .AN(n1312), .B(n1306), .Y(n1305) );
  OAI2BB2X1 U504 ( .B0(n951), .B1(n950), .A0N(n951), .A1N(n950), .Y(n959) );
  NOR2X1 U505 ( .A(n1517), .B(n1516), .Y(n1530) );
  NOR2BX1 U506 ( .AN(n952), .B(n959), .Y(n960) );
  OAI21X1 U507 ( .A0(n223), .A1(n1040), .B0(n1037), .Y(n1043) );
  OA21X2 U508 ( .A0(n209), .A1(n971), .B0(n966), .Y(n974) );
  OAI21X1 U509 ( .A0(n972), .A1(n965), .B0(n209), .Y(n966) );
  AOI32X1 U510 ( .A0(n227), .A1(n1429), .A2(n1412), .B0(n1420), .B1(n1429), 
        .Y(n1431) );
  NOR2X1 U511 ( .A(n227), .B(n1412), .Y(n1420) );
  OAI21X1 U512 ( .A0(n262), .A1(n1007), .B0(n1003), .Y(n1005) );
  AOI22X1 U513 ( .A0(n806), .A1(n805), .B0(n804), .B1(n803), .Y(n810) );
  AOI31X1 U514 ( .A0(n790), .A1(n789), .A2(n2156), .B0(n788), .Y(n806) );
  OAI21X1 U515 ( .A0(n227), .A1(n1062), .B0(n1069), .Y(n1064) );
  AOI21X1 U516 ( .A0(n1593), .A1(n1592), .B0(n1595), .Y(n1610) );
  NOR2X1 U517 ( .A(n1039), .B(n1042), .Y(n1045) );
  OAI21X1 U518 ( .A0(n1038), .A1(n1037), .B0(n1036), .Y(n1042) );
  OAI21X1 U519 ( .A0(n458), .A1(n459), .B0(n513), .Y(n520) );
  OAI211X1 U520 ( .A0(n1798), .A1(n1081), .B0(n1080), .C0(n1079), .Y(n1094) );
  OAI211X1 U521 ( .A0(n1286), .A1(n1084), .B0(n1076), .C0(work_cntr[19]), .Y(
        n1080) );
  OAI21X1 U522 ( .A0(n277), .A1(read_cntr[1]), .B0(n424), .Y(n617) );
  OAI22X1 U523 ( .A0(n1164), .A1(n1169), .B0(n1163), .B1(n1162), .Y(n1173) );
  OAI21X1 U524 ( .A0(n1157), .A1(n1151), .B0(n1165), .Y(n1163) );
  NOR2BX2 U525 ( .AN(n1055), .B(n1054), .Y(n1065) );
  NOR2X1 U526 ( .A(n1052), .B(n1051), .Y(n1054) );
  OAI21X1 U527 ( .A0(write_addr[7]), .A1(n1965), .B0(n1964), .Y(n2101) );
  OAI21X1 U528 ( .A0(n834), .A1(n833), .B0(n832), .Y(n856) );
  OAI2BB2X1 U529 ( .B0(n410), .B1(n2101), .A0N(n2108), .A1N(n2102), .Y(n583)
         );
  OAI21X1 U530 ( .A0(n1599), .A1(n1610), .B0(n1598), .Y(n1603) );
  OAI21X1 U531 ( .A0(write_addr[18]), .A1(n1962), .B0(n1969), .Y(n2213) );
  OAI21X1 U532 ( .A0(n1382), .A1(n1381), .B0(n1380), .Y(n1385) );
  OAI22X1 U533 ( .A0(n901), .A1(n900), .B0(n909), .B1(n899), .Y(n1986) );
  NAND2X1 U534 ( .A(n728), .B(n718), .Y(n909) );
  AOI22X2 U535 ( .A0(n830), .A1(n829), .B0(n828), .B1(n827), .Y(n839) );
  CLKINVX1 U536 ( .A(n1876), .Y(n1880) );
  AOI22X1 U537 ( .A0(work_cntr[8]), .A1(n1864), .B0(n1863), .B1(n1894), .Y(
        n1876) );
  OAI21X1 U538 ( .A0(n989), .A1(n988), .B0(n987), .Y(n995) );
  OAI21X1 U539 ( .A0(n983), .A1(n982), .B0(n269), .Y(n988) );
  OAI21X1 U540 ( .A0(n1831), .A1(n1835), .B0(n1840), .Y(n1838) );
  AOI21X1 U541 ( .A0(n1550), .A1(n1558), .B0(n1554), .Y(n1562) );
  OAI21X1 U542 ( .A0(n957), .A1(n961), .B0(n956), .Y(n964) );
  OAI21X1 U543 ( .A0(n960), .A1(n955), .B0(n268), .Y(n961) );
  OAI21X1 U544 ( .A0(n1525), .A1(n1532), .B0(n1524), .Y(n1533) );
  AOI221X1 U545 ( .A0(n1526), .A1(n1520), .B0(n1527), .B1(n1520), .C0(n1519), 
        .Y(n1525) );
  OAI2BB1X2 U546 ( .A0N(n632), .A1N(n624), .B0(n623), .Y(n625) );
  OAI21X1 U547 ( .A0(n1250), .A1(n1248), .B0(n1247), .Y(n1277) );
  NOR2BX1 U548 ( .AN(n1800), .B(n1813), .Y(n1807) );
  OAI22X2 U549 ( .A0(n2104), .A1(n1935), .B0(n1934), .B1(n2211), .Y(next_en_si) );
  AOI21X1 U550 ( .A0(n2219), .A1(next_en_si), .B0(n149), .Y(n1939) );
  OAI22X1 U551 ( .A0(n1797), .A1(n1796), .B0(work_cntr[19]), .B1(n1799), .Y(
        n1813) );
  NOR2X1 U552 ( .A(work_cntr[11]), .B(n1808), .Y(n1321) );
  OAI21X2 U553 ( .A0(n1479), .A1(n1474), .B0(n1480), .Y(n1488) );
  OAI21X1 U554 ( .A0(n1465), .A1(n1467), .B0(n1464), .Y(n1474) );
  NOR2X1 U555 ( .A(n254), .B(n1204), .Y(n1202) );
  NOR3BX1 U556 ( .AN(n324), .B(write_cntr[12]), .C(n1203), .Y(n1204) );
  NAND2BX1 U557 ( .AN(next_work_cntr[11]), .B(n1499), .Y(n1459) );
  OAI21X1 U558 ( .A0(n2223), .A1(n258), .B0(n2224), .Y(n1201) );
  AOI21X1 U559 ( .A0(n2225), .A1(N1183), .B0(n2224), .Y(n2239) );
  OAI22X1 U560 ( .A0(n1509), .A1(n1508), .B0(n1507), .B1(n1506), .Y(n1516) );
  NAND2X1 U561 ( .A(n481), .B(n512), .Y(n516) );
  CLKINVX1 U562 ( .A(n1640), .Y(n1639) );
  OAI22X2 U563 ( .A0(n1444), .A1(next_cr_x[5]), .B0(n180), .B1(n2082), .Y(
        n1996) );
  NAND3X1 U564 ( .A(n1996), .B(n2006), .C(n1997), .Y(n1991) );
  AOI2BB2X2 U565 ( .B0(n264), .B1(n895), .A0N(n264), .A1N(n895), .Y(n1640) );
  OAI21X1 U566 ( .A0(n1112), .A1(n1111), .B0(n1110), .Y(n1117) );
  AOI2BB2X2 U567 ( .B0(n1996), .B1(n1995), .A0N(n1996), .A1N(n1995), .Y(n2009)
         );
  AOI2BB2X2 U568 ( .B0(n1101), .B1(n1100), .A0N(n1101), .A1N(n1099), .Y(n1111)
         );
  XOR2X1 U569 ( .A(write_addr[6]), .B(n1963), .Y(n2091) );
  NOR2X1 U570 ( .A(n1442), .B(n849), .Y(n851) );
  AOI2BB2X2 U571 ( .B0(n2119), .B1(n1443), .A0N(n2119), .A1N(n1443), .Y(n849)
         );
  AOI2BB2X2 U572 ( .B0(n1892), .B1(n1898), .A0N(n1892), .A1N(n1891), .Y(n1903)
         );
  NOR2X2 U573 ( .A(N1184), .B(n1403), .Y(n1423) );
  NOR4X1 U574 ( .A(global_cntr[7]), .B(global_cntr[10]), .C(global_cntr[13]), 
        .D(global_cntr[15]), .Y(n928) );
  NOR3X2 U575 ( .A(n640), .B(n641), .C(n679), .Y(n1614) );
  OAI21X1 U576 ( .A0(n1968), .A1(write_addr[8]), .B0(n2115), .Y(n2196) );
  NOR4X2 U577 ( .A(global_cntr[0]), .B(global_cntr[1]), .C(n1283), .D(N1593), 
        .Y(en_photo_num) );
  NAND2X1 U578 ( .A(n433), .B(n435), .Y(h_1[2]) );
  NOR2X1 U579 ( .A(n383), .B(n382), .Y(n435) );
  NAND2X1 U580 ( .A(n1960), .B(write_addr[13]), .Y(n2199) );
  NOR2X1 U581 ( .A(n1898), .B(n1890), .Y(n1904) );
  OAI22X1 U582 ( .A0(n1904), .A1(n1893), .B0(n178), .B1(n1903), .Y(n1907) );
  NOR2X1 U583 ( .A(n1599), .B(n1601), .Y(n1592) );
  NOR2X1 U584 ( .A(N1183), .B(n149), .Y(n1599) );
  NOR2X1 U585 ( .A(n1476), .B(n1467), .Y(n1471) );
  NOR2X1 U586 ( .A(n1302), .B(n1295), .Y(n1290) );
  NOR2BX1 U587 ( .AN(n2195), .B(n417), .Y(n558) );
  NOR2X1 U588 ( .A(n2120), .B(n2121), .Y(n2122) );
  NAND3X1 U589 ( .A(work_cntr[6]), .B(n1383), .C(n898), .Y(n885) );
  NOR2X1 U590 ( .A(n223), .B(n229), .Y(n1383) );
  NOR2X1 U591 ( .A(n226), .B(n931), .Y(N1591) );
  OAI31X1 U592 ( .A0(n938), .A1(n937), .A2(n236), .B0(n1077), .Y(n939) );
  OAI31X1 U593 ( .A0(work_cntr[17]), .A1(n259), .A2(n236), .B0(n933), .Y(n941)
         );
  OAI21X1 U594 ( .A0(curr_time[7]), .A1(n873), .B0(n872), .Y(n875) );
  NOR2BX1 U595 ( .AN(n819), .B(n164), .Y(n829) );
  NAND2X1 U596 ( .A(n829), .B(n2184), .Y(n827) );
  OAI21X1 U597 ( .A0(n1844), .A1(n267), .B0(n1824), .Y(n1841) );
  NOR2X1 U598 ( .A(n1808), .B(n1895), .Y(n1844) );
  OAI21X1 U599 ( .A0(n269), .A1(n984), .B0(n988), .Y(n993) );
  OAI21X1 U600 ( .A0(n1843), .A1(n269), .B0(n1808), .Y(n1352) );
  OAI21X1 U601 ( .A0(n1406), .A1(n1403), .B0(N1184), .Y(n1419) );
  AOI2BB2X2 U602 ( .B0(n1460), .B1(next_work_cntr[16]), .A0N(n1460), .A1N(
        next_work_cntr[16]), .Y(n1472) );
  NOR2BX1 U603 ( .AN(n1466), .B(next_work_cntr[15]), .Y(n1460) );
  NOR2X1 U604 ( .A(n778), .B(n779), .Y(n780) );
  OAI31X1 U605 ( .A0(n779), .A1(n778), .A2(n783), .B0(n777), .Y(n791) );
  OAI211X1 U606 ( .A0(n1577), .A1(n1591), .B0(n1582), .C0(n1578), .Y(n1580) );
  NOR2X1 U607 ( .A(n149), .B(work_cntr[4]), .Y(n1577) );
  OAI21X1 U608 ( .A0(n768), .A1(n767), .B0(n766), .Y(n778) );
  NAND2X1 U609 ( .A(n840), .B(n838), .Y(n833) );
  OAI22X1 U610 ( .A0(n177), .A1(n826), .B0(n825), .B1(n824), .Y(n838) );
  OAI22X1 U611 ( .A0(n1559), .A1(n1558), .B0(n1557), .B1(n1556), .Y(n1568) );
  NOR2X1 U612 ( .A(n268), .B(n893), .Y(n894) );
  NAND2X2 U613 ( .A(n215), .B(n894), .Y(n895) );
  NAND2X1 U614 ( .A(n813), .B(n812), .Y(n816) );
  OAI22X1 U615 ( .A0(n2017), .A1(n798), .B0(n797), .B1(n796), .Y(n812) );
  NAND2X1 U616 ( .A(n763), .B(n755), .Y(n770) );
  OAI31X1 U617 ( .A0(n764), .A1(n763), .A2(n765), .B0(n762), .Y(n784) );
  OAI22X1 U618 ( .A0(n750), .A1(n749), .B0(n756), .B1(n748), .Y(n763) );
  NOR2X1 U619 ( .A(n1778), .B(n1195), .Y(n1200) );
  OAI22X1 U620 ( .A0(n1194), .A1(n1193), .B0(n1192), .B1(n1191), .Y(n1195) );
  OAI22X1 U621 ( .A0(n180), .A1(n2143), .B0(n1444), .B1(n2145), .Y(n775) );
  OAI21X1 U622 ( .A0(n775), .A1(n774), .B0(n773), .Y(n789) );
  AOI21X1 U623 ( .A0(work_cntr[18]), .A1(n1288), .B0(n1795), .Y(n1295) );
  NOR2X1 U624 ( .A(n1286), .B(n1289), .Y(n1795) );
  OAI22X1 U625 ( .A0(n2012), .A1(n2011), .B0(n2013), .B1(n2010), .Y(n2035) );
  OAI21X1 U626 ( .A0(n2001), .A1(n2000), .B0(n1999), .Y(n2013) );
  OAI22X1 U627 ( .A0(n1226), .A1(n1225), .B0(n1230), .B1(n1229), .Y(n1246) );
  OAI22X1 U628 ( .A0(n1983), .A1(n1982), .B0(n1984), .B1(n1981), .Y(n2000) );
  OAI21X1 U629 ( .A0(n912), .A1(n911), .B0(n910), .Y(n1984) );
  OAI21X1 U630 ( .A0(n1898), .A1(n1887), .B0(n1897), .Y(n1890) );
  AOI2BB2X2 U631 ( .B0(work_cntr[6]), .B1(n1885), .A0N(work_cntr[6]), .A1N(
        n1885), .Y(n1898) );
  OAI21X1 U632 ( .A0(n771), .A1(n770), .B0(n769), .Y(n776) );
  AOI211X4 U633 ( .A0(n659), .A1(n1940), .B0(n660), .C0(n1939), .Y(n1942) );
  OAI2BB2X1 U634 ( .B0(n2114), .B1(n2113), .A0N(\DP_OP_436J1_125_1438/n26 ), 
        .A1N(n2112), .Y(n2120) );
  NOR2X1 U635 ( .A(n1375), .B(n1374), .Y(n1387) );
  OAI31X4 U636 ( .A0(n1373), .A1(n1372), .A2(n1371), .B0(n1370), .Y(n1374) );
  OAI31X1 U637 ( .A0(n784), .A1(n783), .A2(n782), .B0(n781), .Y(n787) );
  OAI22X1 U638 ( .A0(work_cntr[4]), .A1(n1172), .B0(n223), .B1(n1171), .Y(
        n1177) );
  NAND2BX1 U639 ( .AN(n1301), .B(n1172), .Y(n1090) );
  NOR2X2 U640 ( .A(N1184), .B(n897), .Y(n1172) );
  NOR3X2 U641 ( .A(n258), .B(n228), .C(n1896), .Y(n898) );
  CLKINVX1 U642 ( .A(n1911), .Y(n1896) );
  OAI21X2 U643 ( .A0(n1896), .A1(n228), .B0(n1895), .Y(n1919) );
  AND3X2 U644 ( .A(si_sel), .B(n1431), .C(n1415), .Y(expand_sel[1]) );
  NAND2X1 U645 ( .A(n1233), .B(n1279), .Y(n1240) );
  AND2X2 U646 ( .A(n1279), .B(write_cntr[6]), .Y(n1257) );
  NOR2X1 U647 ( .A(write_cntr[6]), .B(n1279), .Y(n1255) );
  NOR2X1 U648 ( .A(n1279), .B(n430), .Y(n453) );
  CLKINVX1 U649 ( .A(\next_cr_y[0] ), .Y(n170) );
  NOR2X1 U650 ( .A(n1456), .B(n149), .Y(next_work_cntr[19]) );
  OAI21X1 U651 ( .A0(n1474), .A1(n1480), .B0(n1488), .Y(n1484) );
  OAI21X1 U652 ( .A0(n1065), .A1(n1061), .B0(n227), .Y(n1069) );
  AND2X2 U653 ( .A(n656), .B(global_cntr[3]), .Y(n361) );
  AND2X2 U654 ( .A(n657), .B(global_cntr[2]), .Y(n656) );
  OAI21X1 U655 ( .A0(n1861), .A1(n1870), .B0(n1878), .Y(n1877) );
  OAI22X2 U656 ( .A0(n1848), .A1(n265), .B0(n1847), .B1(n1895), .Y(n1870) );
  OAI2BB2X1 U657 ( .B0(n1458), .B1(next_work_cntr[10]), .A0N(n1458), .A1N(
        next_work_cntr[10]), .Y(n1519) );
  NOR2BX1 U658 ( .AN(n1458), .B(next_work_cntr[10]), .Y(n1499) );
  NOR2X2 U659 ( .A(n149), .B(n1691), .Y(next_work_cntr[10]) );
  OAI21X1 U660 ( .A0(n2026), .A1(n163), .B0(n2024), .Y(n2031) );
  NOR3BX1 U661 ( .AN(n163), .B(n2019), .C(n2021), .Y(n2027) );
  NAND3X1 U662 ( .A(n163), .B(n2006), .C(n2017), .Y(n2008) );
  OAI2BB2X1 U663 ( .B0(curr_time[4]), .B1(s_1[3]), .A0N(curr_time[4]), .A1N(
        s_1[3]), .Y(n878) );
  CLKINVX1 U664 ( .A(curr_time[2]), .Y(n658) );
  OAI21X1 U665 ( .A0(n1889), .A1(n1888), .B0(n1887), .Y(n1892) );
  OAI21X2 U666 ( .A0(n1865), .A1(n261), .B0(n1864), .Y(n1888) );
  NOR2X1 U667 ( .A(n2002), .B(n2083), .Y(n2018) );
  CLKINVX1 U668 ( .A(n2017), .Y(n2002) );
  NOR2X2 U669 ( .A(n278), .B(n171), .Y(n2127) );
  NAND2X1 U670 ( .A(cr_read_cntr[5]), .B(n917), .Y(n921) );
  OAI21X1 U671 ( .A0(n914), .A1(n286), .B0(n913), .Y(n917) );
  OAI21X1 U672 ( .A0(n1851), .A1(n1850), .B0(n1849), .Y(n1855) );
  OAI22X1 U673 ( .A0(n1839), .A1(n1850), .B0(n1838), .B1(n1837), .Y(n1852) );
  OAI2BB2X2 U674 ( .B0(work_cntr[12]), .B1(n1824), .A0N(work_cntr[12]), .A1N(
        n1824), .Y(n1850) );
  NOR2X1 U675 ( .A(n1523), .B(n1522), .Y(n1513) );
  NAND2X1 U676 ( .A(n1511), .B(n1510), .Y(n1522) );
  OA21X1 U677 ( .A0(global_cntr[8]), .A1(n365), .B0(n673), .Y(n650) );
  NOR2X2 U678 ( .A(n673), .B(n233), .Y(n648) );
  AOI211X1 U679 ( .A0(n233), .A1(n673), .B0(n648), .C0(n375), .Y(n649) );
  NAND2X1 U680 ( .A(n365), .B(global_cntr[8]), .Y(n673) );
  CLKINVX1 U681 ( .A(n730), .Y(n712) );
  CLKINVX1 U682 ( .A(n1448), .Y(n730) );
  NAND2X1 U683 ( .A(work_cntr[19]), .B(n935), .Y(n1077) );
  NAND2X1 U684 ( .A(n1207), .B(n1281), .Y(n1210) );
  AOI2BB2X2 U685 ( .B0(next_work_cntr[7]), .B1(n1543), .A0N(next_work_cntr[7]), 
        .A1N(n1543), .Y(n1563) );
  NOR2X1 U686 ( .A(n1543), .B(next_work_cntr[7]), .Y(n1536) );
  OAI21X2 U687 ( .A0(n1545), .A1(n1544), .B0(n1543), .Y(n1567) );
  NAND2X1 U688 ( .A(n1545), .B(n1544), .Y(n1543) );
  OAI21X1 U689 ( .A0(n1106), .A1(n1114), .B0(n1122), .Y(n1119) );
  OAI21X2 U690 ( .A0(n1091), .A1(n268), .B0(n1090), .Y(n1114) );
  OAI21X1 U691 ( .A0(work_cntr[8]), .A1(n888), .B0(n889), .Y(n1711) );
  NOR2X1 U692 ( .A(n265), .B(n889), .Y(n890) );
  OAI2BB2X2 U693 ( .B0(n265), .B1(n889), .A0N(n265), .A1N(n889), .Y(n1698) );
  NAND2X1 U694 ( .A(work_cntr[8]), .B(n888), .Y(n889) );
  AOI2BB2X2 U695 ( .B0(n1542), .B1(n1396), .A0N(n1542), .A1N(n1396), .Y(n1404)
         );
  NOR2X1 U696 ( .A(n1397), .B(n1396), .Y(n1402) );
  OAI21X2 U697 ( .A0(n1390), .A1(n1389), .B0(n1388), .Y(n1396) );
  NAND2X1 U698 ( .A(curr_photo_size[0]), .B(curr_photo_size[1]), .Y(n1933) );
  NOR2X1 U699 ( .A(n1915), .B(n1908), .Y(n1913) );
  AOI21X1 U700 ( .A0(n1915), .A1(n1914), .B0(n1913), .Y(n1918) );
  OAI22X2 U701 ( .A0(work_cntr[4]), .A1(n1894), .B0(n223), .B1(n1895), .Y(
        n1915) );
  NOR2X1 U702 ( .A(n149), .B(n1542), .Y(n1569) );
  CLKINVX1 U703 ( .A(n1397), .Y(n1542) );
  OAI21X1 U704 ( .A0(n1153), .A1(n229), .B0(n1152), .Y(n1166) );
  NOR2X1 U705 ( .A(n1152), .B(work_cntr[6]), .Y(n1140) );
  OAI2BB2X2 U706 ( .B0(work_cntr[6]), .B1(n1152), .A0N(work_cntr[6]), .A1N(
        n1152), .Y(n1169) );
  NAND2X1 U707 ( .A(n1791), .B(n1172), .Y(n1152) );
  AOI2BB2X2 U708 ( .B0(next_work_cntr[12]), .B1(n1459), .A0N(
        next_work_cntr[12]), .A1N(n1459), .Y(n1501) );
  NOR2X1 U709 ( .A(next_work_cntr[12]), .B(n1459), .Y(n1486) );
  NOR2X2 U710 ( .A(n149), .B(n1671), .Y(next_work_cntr[12]) );
  CLKINVX1 U711 ( .A(n1447), .Y(n708) );
  OAI211X4 U712 ( .A0(write_cntr[11]), .A1(n705), .B0(n704), .C0(n220), .Y(
        n1447) );
  NAND3X1 U713 ( .A(n1253), .B(n1249), .C(n1261), .Y(n1250) );
  AOI2BB2X2 U714 ( .B0(n1239), .B1(n1238), .A0N(n1239), .A1N(n1238), .Y(n1261)
         );
  NOR2X2 U715 ( .A(work_cntr[16]), .B(n1790), .Y(n1287) );
  NOR2X1 U716 ( .A(n1790), .B(n1895), .Y(n1803) );
  NAND2X1 U717 ( .A(n1809), .B(n264), .Y(n1790) );
  OAI31X4 U718 ( .A0(n1591), .A1(n1590), .A2(n1589), .B0(n1588), .Y(n1595) );
  OAI31X1 U719 ( .A0(n1591), .A1(n1582), .A2(n1581), .B0(n1580), .Y(n1584) );
  NOR2X2 U720 ( .A(n1569), .B(n1565), .Y(n1591) );
  NOR3X2 U721 ( .A(n253), .B(n719), .C(n844), .Y(n724) );
  NOR2X1 U722 ( .A(n837), .B(n844), .Y(n822) );
  NAND2X1 U723 ( .A(write_cntr[1]), .B(write_cntr[0]), .Y(n844) );
  OAI21X2 U724 ( .A0(n1321), .A1(n209), .B0(n1320), .Y(n1337) );
  NAND2X1 U725 ( .A(n1321), .B(n209), .Y(n1320) );
  OAI21X1 U726 ( .A0(n1045), .A1(n1044), .B0(n228), .Y(n1049) );
  OAI21X1 U727 ( .A0(n228), .A1(n1050), .B0(n1049), .Y(n1056) );
  NOR3X1 U728 ( .A(n1408), .B(n228), .C(n1404), .Y(n1406) );
  NAND2X1 U729 ( .A(n222), .B(n236), .Y(n1286) );
  NAND2X1 U730 ( .A(n1287), .B(n222), .Y(n1288) );
  OAI21X2 U731 ( .A0(n1287), .A1(n222), .B0(n1288), .Y(n1298) );
  INVXL U732 ( .A(n1470), .Y(n172) );
  CLKINVX1 U733 ( .A(n172), .Y(n173) );
  NOR2X2 U734 ( .A(n149), .B(n1698), .Y(next_work_cntr[9]) );
  OAI21X1 U735 ( .A0(n1698), .A1(n1697), .B0(n1702), .Y(n1706) );
  NOR2X1 U736 ( .A(n149), .B(n1738), .Y(next_work_cntr[5]) );
  OAI21X1 U737 ( .A0(n1738), .A1(n1737), .B0(n1742), .Y(n1746) );
  OAI21X2 U738 ( .A0(work_cntr[5]), .A1(n887), .B0(n886), .Y(n1738) );
  OAI21X1 U739 ( .A0(n1449), .A1(n735), .B0(n734), .Y(n742) );
  NAND2X1 U740 ( .A(n701), .B(n220), .Y(n1449) );
  CLKINVX1 U741 ( .A(n1778), .Y(n1783) );
  OAI21X2 U742 ( .A0(n847), .A1(n271), .B0(n846), .Y(n1442) );
  NAND2X1 U743 ( .A(n220), .B(n837), .Y(n847) );
  CLKINVX1 U744 ( .A(n1951), .Y(n1947) );
  AOI32X1 U745 ( .A0(cr_read_cntr[6]), .A1(n1952), .A2(cr_read_cntr[7]), .B0(
        n1951), .B1(n1952), .Y(n1953) );
  NAND2X1 U746 ( .A(n1938), .B(next_en_si), .Y(n1951) );
  CLKINVX1 U747 ( .A(n530), .Y(n174) );
  NOR2X1 U748 ( .A(n1563), .B(n1571), .Y(n1558) );
  NAND2X1 U749 ( .A(n1549), .B(n1553), .Y(n1571) );
  CLKINVX1 U750 ( .A(n1378), .Y(n175) );
  AOI2BB2X2 U751 ( .B0(work_cntr[13]), .B1(n1811), .A0N(work_cntr[13]), .A1N(
        n1811), .Y(n1835) );
  NOR2X2 U752 ( .A(n149), .B(n1678), .Y(next_work_cntr[11]) );
  OAI2BB2X2 U753 ( .B0(n267), .B1(n891), .A0N(n267), .A1N(n891), .Y(n1678) );
  OAI211X4 U754 ( .A0(write_cntr[2]), .A1(n822), .B0(n220), .C0(n821), .Y(
        n1443) );
  NAND2X1 U755 ( .A(write_cntr[2]), .B(n822), .Y(n821) );
  CLKINVX1 U756 ( .A(n527), .Y(n176) );
  NOR2X2 U757 ( .A(n1418), .B(n2241), .Y(expand_sel[2]) );
  NOR3BX1 U758 ( .AN(n1369), .B(n1365), .C(n1366), .Y(n1360) );
  NOR2X1 U759 ( .A(n1358), .B(n1366), .Y(n1349) );
  NAND2X1 U760 ( .A(n1347), .B(n1346), .Y(n1366) );
  OAI22X1 U761 ( .A0(n1446), .A1(n2138), .B0(n904), .B1(n2140), .Y(n768) );
  OAI22X2 U762 ( .A0(n904), .A1(n2087), .B0(n1446), .B1(next_cr_x[6]), .Y(
        n1977) );
  CLKINVX1 U763 ( .A(n1446), .Y(n904) );
  CLKINVX1 U764 ( .A(n1902), .Y(n178) );
  OAI21X2 U765 ( .A0(n1291), .A1(n1292), .B0(n1304), .Y(n1314) );
  CLKINVX1 U766 ( .A(n2055), .Y(n2077) );
  NAND2X1 U767 ( .A(n2038), .B(n2037), .Y(n2055) );
  CLKINVX1 U768 ( .A(\DP_OP_166J1_126_2191/I3 ), .Y(n179) );
  OAI2BB2X1 U769 ( .B0(n2166), .B1(n2165), .A0N(n2166), .A1N(n2164), .Y(n2171)
         );
  CLKINVX1 U770 ( .A(n2164), .Y(n2163) );
  NOR2X2 U771 ( .A(n795), .B(n800), .Y(n2164) );
  NOR2X2 U772 ( .A(n149), .B(n1633), .Y(next_work_cntr[16]) );
  OA21X2 U773 ( .A0(n1633), .A1(n1634), .B0(n1632), .Y(n1644) );
  OAI21X1 U774 ( .A0(n1635), .A1(n1631), .B0(n1633), .Y(n1632) );
  OAI21X2 U775 ( .A0(work_cntr[16]), .A1(n896), .B0(n1627), .Y(n1633) );
  OAI31X4 U776 ( .A0(n851), .A1(n2040), .A2(n852), .B0(n856), .Y(n2124) );
  NAND2BX1 U777 ( .AN(n2040), .B(n2039), .Y(n2041) );
  AOI22X2 U778 ( .A0(n836), .A1(n835), .B0(n839), .B1(n843), .Y(n2040) );
  OAI22X1 U779 ( .A0(n1766), .A1(n1197), .B0(n2235), .B1(n1196), .Y(n1199) );
  CLKINVX1 U780 ( .A(n1766), .Y(n2235) );
  AOI2BB1X2 U781 ( .A0N(write_cntr[6]), .A1N(n725), .B0(n726), .Y(n1997) );
  NAND3X1 U782 ( .A(write_cntr[6]), .B(n1239), .C(n1234), .Y(n1233) );
  NOR2X1 U783 ( .A(N1182), .B(n149), .Y(n1606) );
  OA22XL U784 ( .A0(n837), .A1(n717), .B0(n245), .B1(n847), .Y(n1975) );
  INVX3 U785 ( .A(n1975), .Y(n180) );
  CLKINVX1 U786 ( .A(n180), .Y(n1444) );
  INVX4 U787 ( .A(n48), .Y(n334) );
  NAND2X1 U788 ( .A(work_cntr[10]), .B(n890), .Y(n891) );
  OAI21X2 U789 ( .A0(work_cntr[10]), .A1(n890), .B0(n891), .Y(n1691) );
  NAND2X1 U790 ( .A(n809), .B(n2021), .Y(n813) );
  NOR2X1 U791 ( .A(n2078), .B(n2021), .Y(n2020) );
  OAI211X4 U792 ( .A0(write_cntr[4]), .A1(n807), .B0(n220), .C0(n720), .Y(
        n2021) );
  OAI22X1 U793 ( .A0(n908), .A1(n2135), .B0(n737), .B1(n2136), .Y(n750) );
  NOR2X1 U794 ( .A(n905), .B(n908), .Y(n713) );
  INVX3 U795 ( .A(n737), .Y(n908) );
  NOR2XL U796 ( .A(n257), .B(n1189), .Y(n897) );
  AOI2BB2X4 U797 ( .B0(n257), .B1(n1189), .A0N(n257), .A1N(n1189), .Y(n1766)
         );
  OAI21X1 U798 ( .A0(n1054), .A1(n1053), .B0(n257), .Y(n1059) );
  INVX16 U799 ( .A(n4), .Y(cr_a[2]) );
  INVX16 U800 ( .A(n2), .Y(cr_a[0]) );
  INVX16 U801 ( .A(n3), .Y(cr_a[1]) );
  CLKINVX1 U802 ( .A(n2250), .Y(n184) );
  INVX16 U803 ( .A(n184), .Y(cr_a[3]) );
  CLKINVX1 U804 ( .A(n2249), .Y(n186) );
  INVX16 U805 ( .A(n186), .Y(cr_a[4]) );
  CLKINVX1 U806 ( .A(n2248), .Y(n188) );
  INVX16 U807 ( .A(n188), .Y(cr_a[5]) );
  CLKINVX1 U808 ( .A(n2247), .Y(n190) );
  INVX16 U809 ( .A(n190), .Y(cr_a[6]) );
  CLKINVX1 U810 ( .A(n2246), .Y(n192) );
  INVX16 U811 ( .A(n192), .Y(cr_a[7]) );
  INVX16 U812 ( .A(n5), .Y(cr_a[8]) );
  INVX3 U813 ( .A(n594), .Y(n616) );
  OR2X2 U814 ( .A(n620), .B(read_cntr[0]), .Y(n594) );
  AOI211X1 U815 ( .A0(n235), .A1(n704), .B0(n703), .C0(n149), .Y(n1448) );
  NOR2X2 U816 ( .A(n149), .B(n1652), .Y(next_work_cntr[14]) );
  NOR2X2 U817 ( .A(n149), .B(n1639), .Y(next_work_cntr[15]) );
  NOR2X2 U818 ( .A(n149), .B(n1618), .Y(next_work_cntr[17]) );
  NOR2X1 U819 ( .A(n149), .B(n1621), .Y(next_work_cntr[18]) );
  BUFX16 U820 ( .A(n2245), .Y(im_wen_n) );
  NAND2X1 U821 ( .A(write_cntr[7]), .B(n1280), .Y(n1235) );
  NAND2X1 U822 ( .A(n2062), .B(n2061), .Y(n2058) );
  OAI2BB2X1 U823 ( .B0(n849), .B1(n848), .A0N(n849), .A1N(n848), .Y(n2061) );
  OAI21X1 U824 ( .A0(n996), .A1(n991), .B0(n265), .Y(n997) );
  NAND2BX1 U825 ( .AN(n996), .B(n998), .Y(n1001) );
  NOR2X1 U826 ( .A(n990), .B(n995), .Y(n996) );
  NOR2BX1 U827 ( .AN(n949), .B(n948), .Y(n954) );
  OAI21X1 U828 ( .A0(n946), .A1(n945), .B0(n944), .Y(n948) );
  NOR2X1 U829 ( .A(n2205), .B(n2204), .Y(n2206) );
  OAI21X1 U830 ( .A0(n1221), .A1(n1235), .B0(n1220), .Y(n1222) );
  NOR2X2 U831 ( .A(n1215), .B(n1221), .Y(n1239) );
  NOR2X1 U832 ( .A(write_cntr[8]), .B(n1281), .Y(n1221) );
  NOR2X1 U833 ( .A(n1960), .B(write_addr[13]), .Y(n2200) );
  NOR2X1 U834 ( .A(n1959), .B(n275), .Y(n1960) );
  NAND2X1 U835 ( .A(work_cntr[12]), .B(n892), .Y(n893) );
  OAI21X2 U836 ( .A0(work_cntr[12]), .A1(n892), .B0(n893), .Y(n1671) );
  NOR2X1 U837 ( .A(n267), .B(n891), .Y(n892) );
  NOR2X1 U838 ( .A(n513), .B(curr_time[1]), .Y(n502) );
  NAND2X1 U839 ( .A(n457), .B(n456), .Y(n513) );
  NAND2X1 U840 ( .A(n786), .B(n2004), .Y(n790) );
  CLKINVX1 U841 ( .A(n1997), .Y(n2004) );
  NOR2X1 U842 ( .A(n2066), .B(n238), .Y(n2080) );
  NAND2X1 U843 ( .A(write_addr[2]), .B(write_addr[1]), .Y(n2066) );
  NOR2BX1 U844 ( .AN(n1779), .B(n1777), .Y(n1789) );
  NOR2X1 U845 ( .A(n1775), .B(n1774), .Y(n1777) );
  NOR2X1 U846 ( .A(n1791), .B(n1383), .Y(n1397) );
  NOR2X2 U847 ( .A(work_cntr[4]), .B(work_cntr[5]), .Y(n1791) );
  NAND2BX1 U848 ( .AN(n1394), .B(n1391), .Y(n1401) );
  NOR2X1 U849 ( .A(n1384), .B(n1385), .Y(n1394) );
  NOR2X1 U850 ( .A(n235), .B(n704), .Y(n703) );
  NAND2X1 U851 ( .A(write_cntr[11]), .B(n705), .Y(n704) );
  NAND2X1 U852 ( .A(n195), .B(n196), .Y(n1547) );
  NAND2XL U853 ( .A(n1535), .B(n1534), .Y(n195) );
  NOR2X1 U854 ( .A(n1518), .B(n1530), .Y(n1535) );
  NOR2BX1 U855 ( .AN(n1537), .B(n1533), .Y(n1534) );
  NAND2BX1 U856 ( .AN(n1398), .B(n223), .Y(n1405) );
  OAI31X4 U857 ( .A0(n1395), .A1(n1394), .A2(n1393), .B0(n1392), .Y(n1398) );
  NOR2X1 U858 ( .A(n223), .B(n1457), .Y(n887) );
  NAND2X1 U859 ( .A(n1803), .B(n260), .Y(n1802) );
  OAI21X1 U860 ( .A0(n1830), .A1(n1829), .B0(n1828), .Y(n1834) );
  OAI2BB2X1 U861 ( .B0(curr_time[20]), .B1(h_1[3]), .A0N(curr_time[20]), .A1N(
        h_1[3]), .Y(n864) );
  OAI2BB2X2 U862 ( .B0(n1179), .B1(n1178), .A0N(n1179), .A1N(n1177), .Y(n1188)
         );
  OAI21X1 U863 ( .A0(n1167), .A1(n1166), .B0(n1180), .Y(n1179) );
  OAI21X1 U864 ( .A0(n1004), .A1(n1003), .B0(n1002), .Y(n1012) );
  OAI21X1 U865 ( .A0(n152), .A1(n1742), .B0(n1741), .Y(n1749) );
  OAI22X1 U866 ( .A0(n1859), .A1(n1867), .B0(n1858), .B1(n1857), .Y(n1869) );
  OAI21X1 U867 ( .A0(n1842), .A1(n1841), .B0(n1856), .Y(n1858) );
  NOR2X1 U868 ( .A(n981), .B(n978), .Y(n983) );
  OAI21X1 U869 ( .A0(n974), .A1(n977), .B0(n973), .Y(n981) );
  NAND2X1 U870 ( .A(n197), .B(n198), .Y(n2043) );
  INVXL U871 ( .A(n2059), .Y(n199) );
  INVXL U872 ( .A(n2050), .Y(n200) );
  NAND2XL U873 ( .A(n2050), .B(n2059), .Y(n197) );
  NAND2X1 U874 ( .A(n199), .B(n200), .Y(n198) );
  OAI22X2 U875 ( .A0(write_cntr[0]), .A1(n837), .B0(n272), .B1(n847), .Y(n2050) );
  OAI211X1 U876 ( .A0(n1924), .A1(n1925), .B0(n1923), .C0(n1922), .Y(n1929) );
  NOR2X1 U877 ( .A(n2129), .B(n2128), .Y(n2174) );
  OAI21X1 U878 ( .A0(n2126), .A1(write_addr[10]), .B0(n2125), .Y(n2129) );
  OAI21X1 U879 ( .A0(n1257), .A1(n1264), .B0(n1256), .Y(n1258) );
  NOR2X1 U880 ( .A(n155), .B(n253), .Y(n1264) );
  NOR2BX1 U881 ( .AN(n2100), .B(n2099), .Y(n2110) );
  OAI22X1 U882 ( .A0(n2098), .A1(\intadd_3/n1 ), .B0(n2097), .B1(n2096), .Y(
        n2099) );
  NOR2X1 U883 ( .A(n1936), .B(n2211), .Y(n1937) );
  AOI211X1 U884 ( .A0(n1275), .A1(n1274), .B0(n1273), .C0(n1272), .Y(n1439) );
  NOR2X1 U885 ( .A(n1501), .B(n1500), .Y(n1515) );
  NOR2X1 U886 ( .A(n711), .B(n712), .Y(n710) );
  NOR3X1 U887 ( .A(n1446), .B(n1447), .C(n908), .Y(n711) );
  CLKINVX1 U888 ( .A(n1711), .Y(n1707) );
  OAI211X4 U889 ( .A0(write_cntr[9]), .A1(n707), .B0(n220), .C0(n706), .Y(
        n1446) );
  NOR2X1 U890 ( .A(n221), .B(n706), .Y(n705) );
  NAND2X1 U891 ( .A(write_cntr[9]), .B(n707), .Y(n706) );
  NOR2X1 U892 ( .A(n391), .B(n390), .Y(n396) );
  NOR2X1 U893 ( .A(n662), .B(n668), .Y(n664) );
  AOI211X4 U894 ( .A0(n225), .A1(n668), .B0(n372), .C0(n375), .Y(n641) );
  NAND2X1 U895 ( .A(global_cntr[15]), .B(n370), .Y(n668) );
  NOR2BX1 U896 ( .AN(n1081), .B(n1078), .Y(n1082) );
  NOR2X1 U897 ( .A(n1288), .B(n1171), .Y(n1078) );
  NOR2X1 U898 ( .A(n1325), .B(n1319), .Y(n1335) );
  NOR2X1 U899 ( .A(n1308), .B(n1309), .Y(n1325) );
  NOR2X1 U900 ( .A(n240), .B(n1944), .Y(n1949) );
  NAND2X1 U901 ( .A(N686), .B(n631), .Y(n1944) );
  NOR2BX1 U902 ( .AN(n801), .B(n799), .Y(n805) );
  NOR2X1 U903 ( .A(n1099), .B(n1098), .Y(n1109) );
  NOR2X1 U904 ( .A(n2188), .B(n2187), .Y(n2192) );
  NOR2BX1 U905 ( .AN(n1957), .B(n2230), .Y(n1956) );
  NOR2X1 U906 ( .A(work_cntr[12]), .B(n1824), .Y(n1811) );
  NAND2X1 U907 ( .A(n1844), .B(n267), .Y(n1824) );
  NOR2BX1 U908 ( .AN(n1502), .B(n1504), .Y(n1514) );
  NOR2X1 U909 ( .A(next_work_cntr[17]), .B(n1461), .Y(n1462) );
  NAND2BX1 U910 ( .AN(next_work_cntr[16]), .B(n1460), .Y(n1461) );
  OAI21X1 U911 ( .A0(curr_time[15]), .A1(n866), .B0(n865), .Y(n868) );
  OAI21X1 U912 ( .A0(curr_time[23]), .A1(n858), .B0(n857), .Y(n860) );
  NOR2BX1 U913 ( .AN(n1524), .B(n1525), .Y(n1541) );
  AOI2BB2X2 U914 ( .B0(n1521), .B1(next_work_cntr[9]), .A0N(n1521), .A1N(
        next_work_cntr[9]), .Y(n1532) );
  NOR2BX1 U915 ( .AN(n1521), .B(next_work_cntr[9]), .Y(n1458) );
  NOR2BX1 U916 ( .AN(n1536), .B(next_work_cntr[8]), .Y(n1521) );
  NOR2X1 U917 ( .A(n1846), .B(n1171), .Y(n1138) );
  CLKINVX1 U918 ( .A(n1172), .Y(n1171) );
  OAI21X1 U919 ( .A0(n1183), .A1(n1182), .B0(n1181), .Y(n1184) );
  OAI2BB2X1 U920 ( .B0(n1176), .B1(n1175), .A0N(n1176), .A1N(n1174), .Y(n1183)
         );
  NOR2X1 U921 ( .A(n1492), .B(n1493), .Y(n1504) );
  NAND2X1 U922 ( .A(n1493), .B(n1492), .Y(n1502) );
  OAI2BB2X1 U923 ( .B0(n1487), .B1(n1486), .A0N(n1487), .A1N(n1486), .Y(n1493)
         );
  OAI21X1 U924 ( .A0(n1300), .A1(n1299), .B0(n1305), .Y(n1323) );
  NOR3BX1 U925 ( .AN(n1299), .B(n1314), .C(n1303), .Y(n1306) );
  OAI21X1 U926 ( .A0(n1809), .A1(n264), .B0(n1790), .Y(n1299) );
  NAND2BX1 U927 ( .AN(n744), .B(n743), .Y(n746) );
  NOR2X1 U928 ( .A(N1182), .B(n1073), .Y(n1066) );
  OAI21X1 U929 ( .A0(n1055), .A1(n257), .B0(n1059), .Y(n1073) );
  OAI21X1 U930 ( .A0(n919), .A1(n918), .B0(n108), .Y(n922) );
  OAI2BB2X1 U931 ( .B0(n2042), .B1(n2041), .A0N(n2042), .A1N(n2041), .Y(n2060)
         );
  OAI22X1 U932 ( .A0(n1990), .A1(n1989), .B0(n1998), .B1(n1988), .Y(n2015) );
  OAI21X1 U933 ( .A0(n1987), .A1(n1986), .B0(n1985), .Y(n1998) );
  AOI211X4 U934 ( .A0(n2163), .A1(n2162), .B0(n2161), .C0(n2160), .Y(n2169) );
  OAI21X1 U935 ( .A0(n2156), .A1(n2155), .B0(n2154), .Y(n2162) );
  OAI21X1 U936 ( .A0(curr_time[18]), .A1(n514), .B0(n442), .Y(n496) );
  OAI21X1 U937 ( .A0(n439), .A1(n444), .B0(n440), .Y(n514) );
  OAI21X1 U938 ( .A0(n941), .A1(n943), .B0(n942), .Y(n949) );
  NOR2BX1 U939 ( .AN(n942), .B(n943), .Y(n947) );
  OAI21X1 U940 ( .A0(n236), .A1(n936), .B0(n1077), .Y(n943) );
  OAI31X4 U941 ( .A0(n1728), .A1(n1727), .A2(n1726), .B0(n1725), .Y(n1735) );
  OAI21X1 U942 ( .A0(n1718), .A1(n1717), .B0(n1722), .Y(n1726) );
  OAI31X4 U943 ( .A0(n1668), .A1(n1667), .A2(n1666), .B0(n1665), .Y(n1675) );
  OAI21X1 U944 ( .A0(n1658), .A1(n1657), .B0(n1662), .Y(n1666) );
  OAI31X4 U945 ( .A0(n1649), .A1(n1648), .A2(n1647), .B0(n1646), .Y(n1655) );
  OAI21X1 U946 ( .A0(n1639), .A1(n1638), .B0(n1643), .Y(n1647) );
  OAI21X1 U947 ( .A0(n268), .A1(n962), .B0(n961), .Y(n968) );
  OAI21X1 U948 ( .A0(n232), .A1(n2194), .B0(n2186), .Y(n2193) );
  OAI21X1 U949 ( .A0(n2184), .A1(n2183), .B0(n2182), .Y(n2194) );
  OAI31X4 U950 ( .A0(n1688), .A1(n1687), .A2(n1686), .B0(n1685), .Y(n1695) );
  OAI21X1 U951 ( .A0(n1678), .A1(n1677), .B0(n1682), .Y(n1686) );
  OAI21X1 U952 ( .A0(n2235), .A1(n1773), .B0(n1772), .Y(n1782) );
  OAI21X1 U953 ( .A0(n1958), .A1(write_addr[11]), .B0(n1959), .Y(n2197) );
  NAND2X1 U954 ( .A(n1958), .B(write_addr[11]), .Y(n1959) );
  NOR2BX1 U955 ( .AN(n1276), .B(n1263), .Y(n1275) );
  OAI22X1 U956 ( .A0(n1253), .A1(n1252), .B0(n1251), .B1(n1250), .Y(n1276) );
  INVX3 U957 ( .A(n2190), .Y(n659) );
  OAI21X1 U958 ( .A0(n2190), .A1(n2067), .B0(n405), .Y(n606) );
  OAI22X1 U959 ( .A0(n2190), .A1(n2117), .B0(n2211), .B1(n412), .Y(n574) );
  NAND3X2 U960 ( .A(n697), .B(n2219), .C(n696), .Y(n2190) );
  OAI21X1 U961 ( .A0(n740), .A1(n739), .B0(n738), .Y(n758) );
  NOR2BX1 U962 ( .AN(n740), .B(n737), .Y(n744) );
  OAI22X1 U963 ( .A0(n2134), .A1(n708), .B0(n219), .B1(n1447), .Y(n740) );
  OAI22X1 U964 ( .A0(n1209), .A1(n1208), .B0(n1217), .B1(n1216), .Y(n1232) );
  AOI221X4 U965 ( .A0(n1341), .A1(n1339), .B0(n1350), .B1(n1339), .C0(n1340), 
        .Y(n1351) );
  AOI2BB2X2 U966 ( .B0(n1338), .B1(n1337), .A0N(n1338), .A1N(n1337), .Y(n1350)
         );
  NOR3X2 U967 ( .A(n837), .B(n719), .C(n844), .Y(n722) );
  NOR2X4 U968 ( .A(n1937), .B(n1938), .Y(n837) );
  MXI2X2 U969 ( .A(n437), .B(n444), .S0(n441), .Y(n515) );
  NOR2X1 U970 ( .A(n443), .B(curr_time[18]), .Y(n444) );
  XOR2X1 U971 ( .A(n465), .B(curr_time[12]), .Y(n871) );
  NAND2X1 U972 ( .A(n385), .B(n467), .Y(n465) );
  NOR2X1 U973 ( .A(n1585), .B(n1584), .Y(n1594) );
  AOI2BB2X2 U974 ( .B0(n1532), .B1(n1531), .A0N(n1532), .A1N(n1531), .Y(n1550)
         );
  OAI31X4 U975 ( .A0(n1530), .A1(n1529), .A2(n1533), .B0(n1528), .Y(n1531) );
  MXI2X2 U976 ( .A(n880), .B(curr_time[3]), .S0(n879), .Y(n881) );
  AND2X2 U977 ( .A(n394), .B(n396), .Y(n879) );
  CLKINVX1 U978 ( .A(n2136), .Y(n2135) );
  NAND2X1 U979 ( .A(n736), .B(n742), .Y(n2136) );
  OAI21X1 U980 ( .A0(n1862), .A1(n262), .B0(n1846), .Y(n1363) );
  NOR2X2 U981 ( .A(work_cntr[9]), .B(n1846), .Y(n1843) );
  NAND2X1 U982 ( .A(n1862), .B(n262), .Y(n1846) );
  OAI21X1 U983 ( .A0(n2141), .A1(n2140), .B0(n2139), .Y(n2147) );
  CLKINVX1 U984 ( .A(n2140), .Y(n2138) );
  NAND2X1 U985 ( .A(n1843), .B(n269), .Y(n1808) );
  AOI22X1 U986 ( .A0(n1575), .A1(n1574), .B0(n1573), .B1(n1580), .Y(n1576) );
  ADDFX2 U987 ( .A(n1563), .B(n1562), .CI(n1566), .CO(n1574), .S(n1573) );
  CLKINVX1 U988 ( .A(n635), .Y(n696) );
  NAND2X1 U989 ( .A(n635), .B(next_state[1]), .Y(n2045) );
  NOR4X1 U990 ( .A(n635), .B(n2220), .C(n2219), .D(n2218), .Y(n2221) );
  NOR2X2 U991 ( .A(n689), .B(n376), .Y(n635) );
  BUFX4 U992 ( .A(n634), .Y(n337) );
  NOR2XL U993 ( .A(en_so), .B(n48), .Y(n634) );
  NAND2BX1 U994 ( .AN(n1333), .B(n1326), .Y(n1341) );
  NOR2X1 U995 ( .A(n1333), .B(n1332), .Y(n1334) );
  NOR2X1 U996 ( .A(n1317), .B(n1318), .Y(n1333) );
  CLKINVX1 U997 ( .A(n2172), .Y(n2184) );
  OAI22X1 U998 ( .A0(n1445), .A1(n2184), .B0(n177), .B1(n2172), .Y(n836) );
  OAI21X1 U999 ( .A0(n1955), .A1(n916), .B0(n915), .Y(n920) );
  NOR2X2 U1000 ( .A(cr_read_cntr[8]), .B(n287), .Y(n1955) );
  AOI21X2 U1001 ( .A0(n1947), .A1(n1946), .B0(n1945), .Y(n1952) );
  OAI21X1 U1002 ( .A0(n1943), .A1(n1951), .B0(n1942), .Y(n1945) );
  NAND2X1 U1003 ( .A(n201), .B(n202), .Y(n1228) );
  CLKINVX1 U1004 ( .A(n1214), .Y(n203) );
  NAND2XL U1005 ( .A(n113), .B(n1214), .Y(n201) );
  NAND2X1 U1006 ( .A(n203), .B(write_cntr[10]), .Y(n202) );
  OAI21X1 U1007 ( .A0(n1213), .A1(n1215), .B0(n1212), .Y(n1214) );
  OAI2BB2X1 U1008 ( .B0(n1228), .B1(n1227), .A0N(n1228), .A1N(n1227), .Y(n1243) );
  NAND3X1 U1009 ( .A(n1226), .B(n1228), .C(n1224), .Y(n1229) );
  NOR2BX2 U1010 ( .AN(n1587), .B(n1579), .Y(n1593) );
  NOR2X1 U1011 ( .A(n1577), .B(n1576), .Y(n1579) );
  NAND2X1 U1012 ( .A(n1577), .B(n1576), .Y(n1587) );
  NOR2X2 U1013 ( .A(write_cntr[5]), .B(n1441), .Y(n1268) );
  NOR2X2 U1014 ( .A(n1379), .B(n1377), .Y(n1386) );
  NOR2X1 U1015 ( .A(n1364), .B(n1363), .Y(n1377) );
  CLKINVX1 U1016 ( .A(n1376), .Y(n1379) );
  OAI21X1 U1017 ( .A0(n1123), .A1(n1129), .B0(n1137), .Y(n1136) );
  NOR2X1 U1018 ( .A(work_cntr[10]), .B(n1124), .Y(n1108) );
  NOR2XL U1019 ( .A(n1138), .B(n265), .Y(n205) );
  CLKINVX1 U1020 ( .A(n1124), .Y(n206) );
  NAND2X1 U1021 ( .A(n1138), .B(n265), .Y(n1124) );
  OAI21X1 U1022 ( .A0(n1144), .A1(n204), .B0(n1150), .Y(n1148) );
  OAI2BB2X1 U1023 ( .B0(n162), .B1(n1145), .A0N(n162), .A1N(n204), .Y(n1156)
         );
  NAND2X1 U1024 ( .A(n207), .B(n208), .Y(n1126) );
  CLKINVX1 U1025 ( .A(n1107), .Y(n210) );
  NAND2XL U1026 ( .A(n1107), .B(work_cntr[12]), .Y(n207) );
  NAND2X1 U1027 ( .A(n209), .B(n210), .Y(n208) );
  NAND2X1 U1028 ( .A(n1108), .B(n267), .Y(n1107) );
  OAI21X1 U1029 ( .A0(n1127), .A1(n1126), .B0(n1125), .Y(n1130) );
  OAI22X1 U1030 ( .A0(n1120), .A1(n1126), .B0(n1119), .B1(n1118), .Y(n1128) );
  NOR2XL U1031 ( .A(n1085), .B(n260), .Y(n212) );
  INVXL U1032 ( .A(n1084), .Y(n213) );
  NAND2X1 U1033 ( .A(n260), .B(n1085), .Y(n1084) );
  BUFX2 U1034 ( .A(n1821), .Y(n214) );
  NOR2BX2 U1035 ( .AN(n1212), .B(n1213), .Y(n1223) );
  NOR2X1 U1036 ( .A(n1278), .B(n230), .Y(n1213) );
  OAI22X2 U1037 ( .A0(n1978), .A1(n2107), .B0(n216), .B1(n2092), .Y(n2006) );
  CLKINVX1 U1038 ( .A(n2107), .Y(n2092) );
  NAND2X2 U1039 ( .A(n1985), .B(n1984), .Y(n2107) );
  CLKINVX1 U1040 ( .A(n671), .Y(n375) );
  NOR2X1 U1041 ( .A(work_cntr[7]), .B(n1285), .Y(n1862) );
  OAI2BB2X1 U1042 ( .B0(n2147), .B1(n2146), .A0N(n2147), .A1N(n2145), .Y(n2153) );
  CLKINVX1 U1043 ( .A(n2145), .Y(n2143) );
  NOR2X2 U1044 ( .A(n761), .B(n760), .Y(n2145) );
  NOR2X2 U1045 ( .A(n150), .B(n2211), .Y(n2090) );
  NAND2X4 U1046 ( .A(n220), .B(n2104), .Y(n2211) );
  AOI22X1 U1047 ( .A0(n659), .A1(\intadd_3/SUM[0] ), .B0(n2075), .B1(n2090), 
        .Y(n2233) );
  CLKINVX1 U1048 ( .A(n2090), .Y(n410) );
  OAI2BB2X1 U1049 ( .B0(n2159), .B1(n2158), .A0N(n2159), .A1N(n2157), .Y(n2166) );
  CLKINVX1 U1050 ( .A(n2157), .Y(n2156) );
  OAI31X4 U1051 ( .A0(n794), .A1(n2157), .A2(n793), .B0(n792), .Y(n800) );
  NOR2X2 U1052 ( .A(n785), .B(n787), .Y(n2157) );
  OAI31X1 U1053 ( .A0(n843), .A1(n842), .A2(n2119), .B0(n841), .Y(n852) );
  NOR2X2 U1054 ( .A(n831), .B(n839), .Y(n2119) );
  NOR2X2 U1055 ( .A(n155), .B(n524), .Y(n529) );
  NAND2BX1 U1056 ( .AN(n452), .B(n453), .Y(n524) );
  OAI21X2 U1057 ( .A0(n1795), .A1(n259), .B0(n1429), .Y(n1293) );
  NAND2X2 U1058 ( .A(n1793), .B(n1287), .Y(n1429) );
  NOR2X1 U1059 ( .A(n1477), .B(n1489), .Y(n1479) );
  NOR3X1 U1060 ( .A(n1485), .B(n1489), .C(n1484), .Y(n1490) );
  OAI21X2 U1061 ( .A0(n1473), .A1(n1472), .B0(n1478), .Y(n1489) );
  OAI2BB2X2 U1062 ( .B0(n1354), .B1(n1353), .A0N(n1354), .A1N(n1353), .Y(n1369) );
  OAI21X1 U1063 ( .A0(n1350), .A1(n1345), .B0(n1344), .Y(n1353) );
  NAND2X1 U1064 ( .A(n1999), .B(n1998), .Y(n2095) );
  CLKINVX1 U1065 ( .A(n2086), .Y(n2083) );
  OAI22X1 U1066 ( .A0(n2018), .A1(n2020), .B0(n2017), .B1(n2086), .Y(n2026) );
  OAI21X2 U1067 ( .A0(n2064), .A1(n2086), .B0(n2076), .Y(n2073) );
  NAND2X2 U1068 ( .A(n2014), .B(n2013), .Y(n2086) );
  AOI21X2 U1069 ( .A0(work_cntr[15]), .A1(n1801), .B0(n1803), .Y(n1816) );
  NOR2X1 U1070 ( .A(n1075), .B(work_cntr[15]), .Y(n1085) );
  OAI22X2 U1071 ( .A0(n264), .A1(n1074), .B0(work_cntr[15]), .B1(n1075), .Y(
        n1089) );
  NAND2X1 U1072 ( .A(n1791), .B(n1894), .Y(n1885) );
  INVX3 U1073 ( .A(n1895), .Y(n1894) );
  NOR2X1 U1074 ( .A(n1766), .B(n1758), .Y(n1414) );
  CLKINVX1 U1075 ( .A(n1758), .Y(n1756) );
  NOR2X1 U1076 ( .A(n1758), .B(n1184), .Y(n1187) );
  NOR2X2 U1077 ( .A(n1172), .B(n898), .Y(n1758) );
  ADDFX2 U1078 ( .A(n2078), .B(n2057), .CI(n2056), .CO(n2074), .S(n2054) );
  NOR2BX2 U1079 ( .AN(n2034), .B(n2036), .Y(n2078) );
  NAND2X2 U1080 ( .A(n228), .B(n1896), .Y(n1895) );
  OAI221X4 U1081 ( .A0(n1921), .A1(n1920), .B0(n1919), .B1(n1918), .C0(n1917), 
        .Y(n1925) );
  OA21X1 U1082 ( .A0(n1910), .A1(n1919), .B0(n1909), .Y(n1924) );
  INVX3 U1083 ( .A(n603), .Y(n613) );
  OR2X2 U1084 ( .A(n2228), .B(n2238), .Y(n603) );
  INVX3 U1085 ( .A(n2167), .Y(n2170) );
  CLKINVX1 U1086 ( .A(n2152), .Y(n783) );
  NAND2X2 U1087 ( .A(n772), .B(n776), .Y(n2152) );
  CLKBUFX3 U1088 ( .A(work_cntr[14]), .Y(n215) );
  OAI21X1 U1089 ( .A0(work_cntr[14]), .A1(n951), .B0(n948), .Y(n953) );
  AOI21X1 U1090 ( .A0(n953), .A1(n949), .B0(n215), .Y(n950) );
  AOI21X1 U1091 ( .A0(n215), .A1(n954), .B0(n950), .Y(n957) );
  NOR2X2 U1092 ( .A(n215), .B(n1301), .Y(n1809) );
  NOR2X1 U1093 ( .A(n1090), .B(n215), .Y(n1074) );
  AOI22X2 U1094 ( .A0(n215), .A1(n1810), .B0(n1809), .B1(n1894), .Y(n1825) );
  OAI2BB2X1 U1095 ( .B0(n215), .B1(n1301), .A0N(n215), .A1N(n1301), .Y(n1308)
         );
  OAI21X2 U1096 ( .A0(n215), .A1(n894), .B0(n895), .Y(n1652) );
  NOR2X1 U1097 ( .A(n256), .B(n726), .Y(n217) );
  NOR2XL U1098 ( .A(write_cntr[7]), .B(n727), .Y(n218) );
  NOR2BX1 U1099 ( .AN(n775), .B(n216), .Y(n779) );
  CLKINVX1 U1100 ( .A(n216), .Y(n1978) );
  NAND3X1 U1101 ( .A(n1977), .B(n1996), .C(n216), .Y(n1979) );
  OAI22X1 U1102 ( .A0(n1994), .A1(n2003), .B0(n216), .B1(n2107), .Y(n1995) );
  CLKINVX1 U1103 ( .A(n608), .Y(n355) );
  OR2X4 U1104 ( .A(n620), .B(n277), .Y(n608) );
  CLKINVX1 U1105 ( .A(next_cr_x[6]), .Y(n2087) );
  INVX3 U1106 ( .A(n718), .Y(next_cr_x[6]) );
  CLKINVX1 U1107 ( .A(next_cr_x[5]), .Y(n2082) );
  NAND2X2 U1108 ( .A(n910), .B(n909), .Y(next_cr_x[5]) );
  AOI221X4 U1109 ( .A0(n1413), .A1(N76), .B0(n1426), .B1(n258), .C0(n2241), 
        .Y(expand_sel[0]) );
  CLKAND2X3 U1110 ( .A(n632), .B(n2228), .Y(n610) );
  BUFX4 U1111 ( .A(n359), .Y(n357) );
  INVX4 U1112 ( .A(n338), .Y(n618) );
  BUFX4 U1113 ( .A(\RSOP_434/C2/CONTROL1 ), .Y(n338) );
  AOI221X4 U1114 ( .A0(n149), .A1(n706), .B0(n221), .B1(n706), .C0(n705), .Y(
        n737) );
  OAI31X4 U1115 ( .A0(n722), .A1(n149), .A2(n253), .B0(n721), .Y(n2017) );
  NOR2X1 U1116 ( .A(n149), .B(n1731), .Y(next_work_cntr[6]) );
  NOR2X2 U1117 ( .A(n149), .B(n1718), .Y(next_work_cntr[7]) );
  INVX6 U1118 ( .A(n147), .Y(n360) );
  NAND2X1 U1119 ( .A(global_cntr[2]), .B(n1282), .Y(n1283) );
  NOR2X2 U1120 ( .A(global_cntr[2]), .B(n931), .Y(N1549) );
  NAND3X1 U1121 ( .A(global_cntr[1]), .B(n1282), .C(n279), .Y(n931) );
  NOR2XL U1122 ( .A(n149), .B(n1778), .Y(next_work_cntr[1]) );
  NOR2XL U1123 ( .A(n149), .B(n1756), .Y(next_work_cntr[3]) );
  NOR2XL U1124 ( .A(n149), .B(n2235), .Y(next_work_cntr[2]) );
  NOR2XL U1125 ( .A(n149), .B(n1753), .Y(next_work_cntr[4]) );
  NAND2XL U1126 ( .A(curr_photo[0]), .B(n325), .Y(n423) );
  NOR2XL U1127 ( .A(curr_photo[0]), .B(n2222), .Y(n2220) );
  NOR3XL U1128 ( .A(n635), .B(n2219), .C(n2218), .Y(n2215) );
  NOR2BXL U1129 ( .AN(N687), .B(n2241), .Y(n2250) );
  NOR2BXL U1130 ( .AN(N688), .B(n2241), .Y(n2249) );
  NOR2BXL U1131 ( .AN(N689), .B(n2241), .Y(n2248) );
  NOR2BXL U1132 ( .AN(N690), .B(n2241), .Y(n2247) );
  NOR2BXL U1133 ( .AN(N691), .B(n2241), .Y(n2246) );
  NAND3XL U1134 ( .A(n494), .B(n493), .C(n492), .Y(\C1/Z_3 ) );
  AOI22XL U1135 ( .A0(n529), .A1(n491), .B0(n176), .B1(s_1[3]), .Y(n492) );
  XNOR2XL U1136 ( .A(n489), .B(n488), .Y(n491) );
  INVXL U1137 ( .A(n483), .Y(n486) );
  NAND2XL U1138 ( .A(n516), .B(n506), .Y(n489) );
  AOI22XL U1139 ( .A0(n174), .A1(h_1[3]), .B0(n528), .B1(n463), .Y(n493) );
  XNOR2XL U1140 ( .A(n462), .B(n461), .Y(n463) );
  NAND2XL U1141 ( .A(n520), .B(n500), .Y(n462) );
  XOR2XL U1142 ( .A(n450), .B(n449), .Y(n451) );
  OAI211XL U1143 ( .A0(n448), .A1(n514), .B0(n447), .C0(n446), .Y(n449) );
  NAND2XL U1144 ( .A(n445), .B(n444), .Y(n447) );
  INVXL U1145 ( .A(n443), .Y(n448) );
  NAND2XL U1146 ( .A(n519), .B(n495), .Y(n450) );
  NAND3XL U1147 ( .A(n510), .B(n509), .C(n508), .Y(\C1/Z_2 ) );
  AOI22XL U1148 ( .A0(n174), .A1(h_1[2]), .B0(n528), .B1(n503), .Y(n509) );
  NAND2BXL U1149 ( .AN(n884), .B(n502), .Y(n500) );
  INVXL U1150 ( .A(n884), .Y(n501) );
  NAND2XL U1151 ( .A(n497), .B(n496), .Y(n495) );
  INVXL U1152 ( .A(n440), .Y(n445) );
  NOR4XL U1153 ( .A(n174), .B(n529), .C(n528), .D(n176), .Y(n533) );
  NAND3XL U1154 ( .A(n523), .B(n522), .C(n521), .Y(\C1/Z_0 ) );
  AOI22XL U1155 ( .A0(\m_0[0] ), .A1(n529), .B0(n176), .B1(n520), .Y(n521) );
  INVXL U1156 ( .A(n883), .Y(n455) );
  NAND2XL U1157 ( .A(n460), .B(n397), .Y(n883) );
  NAND2XL U1158 ( .A(n456), .B(n460), .Y(s_1[1]) );
  NAND2XL U1159 ( .A(n881), .B(n658), .Y(n882) );
  NOR2XL U1160 ( .A(curr_time[3]), .B(n879), .Y(n877) );
  INVXL U1161 ( .A(n876), .Y(n392) );
  NAND2XL U1162 ( .A(n878), .B(n880), .Y(n876) );
  INVXL U1163 ( .A(curr_time[3]), .Y(n880) );
  INVXL U1164 ( .A(n396), .Y(n393) );
  INVXL U1165 ( .A(n389), .Y(n390) );
  NOR2XL U1166 ( .A(curr_time[5]), .B(curr_time[6]), .Y(n874) );
  NOR2XL U1167 ( .A(n388), .B(n387), .Y(n391) );
  INVXL U1168 ( .A(curr_time[6]), .Y(n387) );
  NAND2BXL U1169 ( .AN(n875), .B(n386), .Y(n388) );
  INVXL U1170 ( .A(curr_time[4]), .Y(n386) );
  NAND3XL U1171 ( .A(curr_time[7]), .B(curr_time[6]), .C(n873), .Y(n872) );
  INVXL U1172 ( .A(curr_time[5]), .Y(n873) );
  INVXL U1173 ( .A(curr_time[1]), .Y(n458) );
  AOI22XL U1174 ( .A0(n174), .A1(n519), .B0(n528), .B1(\s_0[0] ), .Y(n522) );
  INVXL U1175 ( .A(n490), .Y(n454) );
  OAI211XL U1176 ( .A0(n439), .A1(curr_time[18]), .B0(n443), .C0(curr_time[17]), .Y(n438) );
  INVXL U1177 ( .A(n439), .Y(n441) );
  INVXL U1178 ( .A(n864), .Y(n436) );
  NAND2XL U1179 ( .A(n446), .B(n440), .Y(n437) );
  NAND2XL U1180 ( .A(n443), .B(curr_time[18]), .Y(n446) );
  INVXL U1181 ( .A(n862), .Y(n431) );
  NAND2XL U1182 ( .A(n861), .B(h_1[2]), .Y(n862) );
  NOR2XL U1183 ( .A(h_1[2]), .B(n861), .Y(n432) );
  INVXL U1184 ( .A(n381), .Y(n382) );
  NOR2XL U1185 ( .A(n380), .B(n379), .Y(n383) );
  INVXL U1186 ( .A(curr_time[22]), .Y(n379) );
  NAND2XL U1187 ( .A(n864), .B(n861), .Y(n863) );
  INVXL U1188 ( .A(curr_time[19]), .Y(n861) );
  NAND2BXL U1189 ( .AN(n860), .B(n378), .Y(n380) );
  INVXL U1190 ( .A(curr_time[20]), .Y(n378) );
  NAND3XL U1191 ( .A(curr_time[23]), .B(curr_time[22]), .C(n858), .Y(n857) );
  INVXL U1192 ( .A(curr_time[21]), .Y(n858) );
  AOI22XL U1193 ( .A0(\h_0[0] ), .A1(n518), .B0(n517), .B1(n516), .Y(n523) );
  INVXL U1194 ( .A(n871), .Y(n480) );
  NAND2XL U1195 ( .A(n477), .B(curr_time[10]), .Y(n478) );
  NAND3XL U1196 ( .A(n483), .B(curr_time[9]), .C(n477), .Y(n481) );
  INVXL U1197 ( .A(n487), .Y(n477) );
  NAND2XL U1198 ( .A(n470), .B(n871), .Y(n471) );
  INVXL U1199 ( .A(n476), .Y(n472) );
  INVXL U1200 ( .A(n870), .Y(n473) );
  NAND2XL U1201 ( .A(n498), .B(curr_time[11]), .Y(n469) );
  INVXL U1202 ( .A(n468), .Y(n498) );
  NAND2XL U1203 ( .A(n468), .B(n869), .Y(n470) );
  NAND2XL U1204 ( .A(n474), .B(n476), .Y(n468) );
  NAND2BXL U1205 ( .AN(n871), .B(n869), .Y(n870) );
  INVXL U1206 ( .A(curr_time[11]), .Y(n869) );
  NOR2XL U1207 ( .A(curr_time[13]), .B(curr_time[14]), .Y(n867) );
  NAND3XL U1208 ( .A(n466), .B(curr_time[14]), .C(n384), .Y(n385) );
  NAND2BXL U1209 ( .AN(curr_time[13]), .B(curr_time[15]), .Y(n384) );
  NAND2BXL U1210 ( .AN(n868), .B(n464), .Y(n466) );
  INVXL U1211 ( .A(curr_time[12]), .Y(n464) );
  NAND3XL U1212 ( .A(curr_time[15]), .B(curr_time[14]), .C(n866), .Y(n865) );
  INVXL U1213 ( .A(curr_time[13]), .Y(n866) );
  INVXL U1214 ( .A(n531), .Y(n517) );
  NAND2BXL U1215 ( .AN(n1280), .B(n429), .Y(n430) );
  NOR2XL U1216 ( .A(n1281), .B(n1202), .Y(n429) );
  AND2XL U1217 ( .A(n452), .B(n428), .Y(n490) );
  NAND2BXL U1218 ( .AN(n1439), .B(n427), .Y(n428) );
  INVXL U1219 ( .A(n1438), .Y(n427) );
  INVXL U1220 ( .A(n1276), .Y(n426) );
  INVXL U1221 ( .A(n1271), .Y(n1272) );
  INVXL U1222 ( .A(n1262), .Y(n1274) );
  INVXL U1223 ( .A(n1255), .Y(n1256) );
  INVXL U1224 ( .A(n1441), .Y(n633) );
  NOR2BXL U1225 ( .AN(n1261), .B(n1260), .Y(n1252) );
  NOR2XL U1226 ( .A(n1241), .B(n1240), .Y(n1242) );
  NAND3XL U1227 ( .A(write_cntr[5]), .B(n1234), .C(n1254), .Y(n1249) );
  INVXL U1228 ( .A(n1235), .Y(n1237) );
  INVXL U1229 ( .A(n1229), .Y(n1231) );
  NOR2BXL U1230 ( .AN(n1228), .B(n1227), .Y(n1225) );
  INVXL U1231 ( .A(n1259), .Y(n1234) );
  NAND2BXL U1232 ( .AN(n1280), .B(n256), .Y(n1236) );
  INVXL U1233 ( .A(n1216), .Y(n1218) );
  NAND3XL U1234 ( .A(write_cntr[7]), .B(n1223), .C(n1239), .Y(n1224) );
  INVXL U1235 ( .A(n1220), .Y(n1215) );
  NAND2XL U1236 ( .A(n1281), .B(write_cntr[8]), .Y(n1220) );
  NOR2XL U1237 ( .A(n166), .B(n1210), .Y(n1208) );
  NAND2XL U1238 ( .A(n1213), .B(write_cntr[10]), .Y(n1205) );
  NAND2XL U1239 ( .A(n230), .B(n1278), .Y(n1212) );
  INVXL U1240 ( .A(n1202), .Y(n1278) );
  NAND2XL U1241 ( .A(n922), .B(n923), .Y(n534) );
  MXI2XL U1242 ( .A(cr_read_cntr[4]), .B(n922), .S0(n923), .Y(n537) );
  AND2XL U1243 ( .A(n535), .B(cr_read_cntr[3]), .Y(n538) );
  NAND2XL U1244 ( .A(n920), .B(n921), .Y(n918) );
  NAND2XL U1245 ( .A(cr_read_cntr[6]), .B(n1955), .Y(n915) );
  NOR2XL U1246 ( .A(n286), .B(n914), .Y(n916) );
  NOR2XL U1247 ( .A(n2237), .B(n1416), .Y(n1417) );
  AOI21XL U1248 ( .A0(n1433), .A1(n1429), .B0(n1428), .Y(n1430) );
  NOR3X1 U1249 ( .A(n2239), .B(n2238), .C(n258), .Y(n2242) );
  INVXL U1250 ( .A(n617), .Y(n425) );
  NAND2XL U1251 ( .A(n1937), .B(next_en_si), .Y(n2244) );
  NOR2XL U1252 ( .A(n1941), .B(n401), .Y(n315) );
  NAND2XL U1253 ( .A(n631), .B(n224), .Y(n402) );
  INVXL U1254 ( .A(n1944), .Y(n403) );
  NAND2XL U1255 ( .A(n360), .B(n615), .Y(n422) );
  NAND2XL U1256 ( .A(write_addr[1]), .B(n266), .Y(n404) );
  NOR2XL U1257 ( .A(n1948), .B(n1952), .Y(n311) );
  AOI21XL U1258 ( .A0(n1949), .A1(cr_read_cntr[4]), .B0(cr_read_cntr[5]), .Y(
        n1948) );
  NAND2XL U1259 ( .A(cr_read_cntr[5]), .B(cr_read_cntr[4]), .Y(n1946) );
  NAND3XL U1260 ( .A(cr_read_cntr[5]), .B(cr_read_cntr[4]), .C(n1949), .Y(
        n1950) );
  XOR2XL U1261 ( .A(n1927), .B(n1926), .Y(n1928) );
  NAND3XL U1262 ( .A(n1924), .B(N1183), .C(n227), .Y(n1922) );
  OAI211XL U1263 ( .A0(n1919), .A1(n1916), .B0(n1920), .C0(n1918), .Y(n1917)
         );
  NAND2XL U1264 ( .A(n1919), .B(n1916), .Y(n1921) );
  NAND2BXL U1265 ( .AN(n1920), .B(n1919), .Y(n1909) );
  NAND2BXL U1266 ( .AN(n1914), .B(n1905), .Y(n1908) );
  NOR2XL U1267 ( .A(n1904), .B(n1900), .Y(n1901) );
  NAND2XL U1268 ( .A(n178), .B(n1903), .Y(n1893) );
  NOR2XL U1269 ( .A(work_cntr[4]), .B(n1895), .Y(n1886) );
  INVXL U1270 ( .A(n1888), .Y(n1883) );
  NAND3XL U1271 ( .A(n1889), .B(n1888), .C(n1879), .Y(n1887) );
  NAND3XL U1272 ( .A(n1881), .B(n1880), .C(n1878), .Y(n1879) );
  INVXL U1273 ( .A(n1881), .Y(n1874) );
  INVXL U1274 ( .A(n1871), .Y(n1873) );
  NOR2XL U1275 ( .A(work_cntr[6]), .B(n1885), .Y(n1865) );
  NAND2XL U1276 ( .A(n1862), .B(n1894), .Y(n1864) );
  NAND3XL U1277 ( .A(n1861), .B(n1870), .C(n1866), .Y(n1878) );
  NAND2BXL U1278 ( .AN(n1860), .B(n1867), .Y(n1866) );
  INVXL U1279 ( .A(n1869), .Y(n1861) );
  NAND2XL U1280 ( .A(n1868), .B(n1856), .Y(n1860) );
  NOR2XL U1281 ( .A(n1846), .B(n1895), .Y(n1848) );
  NAND2XL U1282 ( .A(n1843), .B(n1894), .Y(n1845) );
  INVXL U1283 ( .A(n1858), .Y(n1859) );
  NAND3XL U1284 ( .A(n1842), .B(n1841), .C(n1849), .Y(n1856) );
  NAND3XL U1285 ( .A(n1851), .B(n1850), .C(n1840), .Y(n1849) );
  INVXL U1286 ( .A(n1852), .Y(n1842) );
  INVXL U1287 ( .A(n1831), .Y(n1832) );
  INVXL U1288 ( .A(n1834), .Y(n1836) );
  INVXL U1289 ( .A(n1841), .Y(n1854) );
  INVXL U1290 ( .A(n1838), .Y(n1839) );
  NAND3XL U1291 ( .A(n1831), .B(n1835), .C(n1823), .Y(n1840) );
  NAND3XL U1292 ( .A(n1826), .B(n1830), .C(n1827), .Y(n1823) );
  NAND2XL U1293 ( .A(n1822), .B(n214), .Y(n1827) );
  INVXL U1294 ( .A(n1825), .Y(n1830) );
  INVXL U1295 ( .A(n1829), .Y(n1826) );
  NAND2XL U1296 ( .A(n1811), .B(n268), .Y(n1810) );
  OAI2BB2XL U1297 ( .B0(n1807), .B1(n1806), .A0N(n1807), .A1N(n1805), .Y(n1821) );
  INVXL U1298 ( .A(n1805), .Y(n1812) );
  INVXL U1299 ( .A(n1816), .Y(n1822) );
  NAND2XL U1300 ( .A(n1809), .B(n1894), .Y(n1801) );
  AND2XL U1301 ( .A(n1800), .B(n1815), .Y(n1804) );
  NAND2BXL U1302 ( .AN(n1799), .B(n1798), .Y(n1815) );
  NAND2XL U1303 ( .A(n1797), .B(n1796), .Y(n1800) );
  NOR2XL U1304 ( .A(work_cntr[17]), .B(n1802), .Y(n1794) );
  NAND2XL U1305 ( .A(n1787), .B(n1786), .Y(n1788) );
  NAND2XL U1306 ( .A(n1782), .B(n1780), .Y(n1781) );
  INVXL U1307 ( .A(n1784), .Y(n1776) );
  NOR2XL U1308 ( .A(n1783), .B(n1782), .Y(n1774) );
  NAND2XL U1309 ( .A(n1775), .B(n1784), .Y(n1779) );
  NAND2XL U1310 ( .A(n161), .B(n1769), .Y(n1773) );
  NAND2XL U1311 ( .A(n1765), .B(n1764), .Y(n1769) );
  NOR2XL U1312 ( .A(n1766), .B(n1757), .Y(n1763) );
  INVXL U1313 ( .A(n1757), .Y(n1768) );
  NAND2XL U1314 ( .A(n168), .B(n1754), .Y(n1765) );
  NAND2XL U1315 ( .A(n1762), .B(n1756), .Y(n1754) );
  NAND2BXL U1316 ( .AN(n168), .B(n1759), .Y(n1764) );
  NAND2XL U1317 ( .A(n1750), .B(n1752), .Y(n1759) );
  NAND2XL U1318 ( .A(n1749), .B(n1748), .Y(n1752) );
  NAND2XL U1319 ( .A(n1746), .B(n1751), .Y(n1745) );
  NOR2XL U1320 ( .A(n1747), .B(n1746), .Y(n1744) );
  INVXL U1321 ( .A(n1738), .Y(n1739) );
  NAND2XL U1322 ( .A(n1736), .B(n1737), .Y(n1748) );
  NAND2BXL U1323 ( .AN(n1735), .B(n1740), .Y(n1737) );
  NAND2XL U1324 ( .A(n1734), .B(n1733), .Y(n1740) );
  NAND2XL U1325 ( .A(n1735), .B(n1732), .Y(n1736) );
  NAND2XL U1326 ( .A(n152), .B(n1738), .Y(n1732) );
  NAND2XL U1327 ( .A(n159), .B(n1728), .Y(n1733) );
  NAND2XL U1328 ( .A(n1726), .B(n1730), .Y(n1725) );
  NOR2XL U1329 ( .A(n1727), .B(n1726), .Y(n1724) );
  INVXL U1330 ( .A(n1731), .Y(n1727) );
  NAND2BXL U1331 ( .AN(n1715), .B(n1720), .Y(n1717) );
  NAND2XL U1332 ( .A(n1714), .B(n1713), .Y(n1720) );
  NAND2XL U1333 ( .A(n1715), .B(n1712), .Y(n1716) );
  NAND2XL U1334 ( .A(n1723), .B(n1718), .Y(n1712) );
  NAND2XL U1335 ( .A(n158), .B(n1708), .Y(n1713) );
  NAND2XL U1336 ( .A(n1706), .B(n1710), .Y(n1705) );
  NOR2XL U1337 ( .A(n1707), .B(n1706), .Y(n1704) );
  INVXL U1338 ( .A(n1698), .Y(n1699) );
  NAND2BXL U1339 ( .AN(n1695), .B(n1700), .Y(n1697) );
  NAND2XL U1340 ( .A(n1694), .B(n1693), .Y(n1700) );
  NAND2XL U1341 ( .A(n1695), .B(n1692), .Y(n1696) );
  NAND2XL U1342 ( .A(n1703), .B(n1698), .Y(n1692) );
  NAND2XL U1343 ( .A(n157), .B(n1688), .Y(n1693) );
  NAND2XL U1344 ( .A(n1686), .B(n1690), .Y(n1685) );
  NOR2XL U1345 ( .A(n1687), .B(n1686), .Y(n1684) );
  INVXL U1346 ( .A(n1678), .Y(n1679) );
  INVXL U1347 ( .A(n1691), .Y(n1687) );
  NAND2BXL U1348 ( .AN(n1675), .B(n1680), .Y(n1677) );
  NAND2XL U1349 ( .A(n1674), .B(n1673), .Y(n1680) );
  NAND2XL U1350 ( .A(n1675), .B(n1672), .Y(n1676) );
  NAND2XL U1351 ( .A(n1683), .B(n1678), .Y(n1672) );
  NAND2XL U1352 ( .A(n156), .B(n1668), .Y(n1673) );
  NAND2XL U1353 ( .A(n1666), .B(n1670), .Y(n1665) );
  NOR2XL U1354 ( .A(n1667), .B(n1666), .Y(n1664) );
  INVXL U1355 ( .A(n1671), .Y(n1667) );
  NAND2BXL U1356 ( .AN(n1655), .B(n1660), .Y(n1657) );
  NAND2XL U1357 ( .A(n1654), .B(n1653), .Y(n1660) );
  NAND2XL U1358 ( .A(n1650), .B(n1649), .Y(n1653) );
  NAND2XL U1359 ( .A(n1647), .B(n1651), .Y(n1646) );
  NOR2XL U1360 ( .A(n1648), .B(n1647), .Y(n1645) );
  INVXL U1361 ( .A(n1652), .Y(n1648) );
  NAND2BXL U1362 ( .AN(n1636), .B(n1641), .Y(n1638) );
  NAND2BXL U1363 ( .AN(n1631), .B(n1630), .Y(n1634) );
  NOR2XL U1364 ( .A(n1620), .B(n1619), .Y(n1622) );
  NOR2BXL U1365 ( .AN(n1633), .B(n1629), .Y(n1624) );
  INVXL U1366 ( .A(n1618), .Y(n1620) );
  AOI32XL U1367 ( .A0(n153), .A1(si_sel), .A2(n1617), .B0(n1616), .B1(n2241), 
        .Y(n1935) );
  NOR3XL U1368 ( .A(n635), .B(n2219), .C(next_glb_cntr[2]), .Y(n1615) );
  AOI211XL U1369 ( .A0(n1607), .A1(n1606), .B0(n1605), .C0(n1604), .Y(n1608)
         );
  INVXL U1370 ( .A(n1607), .Y(n1600) );
  NAND2BXL U1371 ( .AN(n1595), .B(n1599), .Y(n1598) );
  INVXL U1372 ( .A(n1601), .Y(n1597) );
  INVXL U1373 ( .A(n1592), .Y(n1609) );
  NAND2XL U1374 ( .A(n1587), .B(n1586), .Y(n1590) );
  NAND2XL U1375 ( .A(n1594), .B(n1593), .Y(n1586) );
  AOI211XL U1376 ( .A0(n1585), .A1(n1587), .B0(n1589), .C0(n1579), .Y(n1581)
         );
  INVXL U1377 ( .A(n1578), .Y(n1589) );
  INVXL U1378 ( .A(n1585), .Y(n1583) );
  INVXL U1379 ( .A(n1574), .Y(n1570) );
  INVXL U1380 ( .A(n1571), .Y(n1572) );
  NAND2XL U1381 ( .A(n1567), .B(n1568), .Y(n1566) );
  NOR2XL U1382 ( .A(n1567), .B(n1568), .Y(n1560) );
  OAI211XL U1383 ( .A0(n1555), .A1(n1554), .B0(n1553), .C0(n1552), .Y(n1557)
         );
  INVXL U1384 ( .A(n1567), .Y(n1551) );
  INVXL U1385 ( .A(n1563), .Y(n1555) );
  NAND2XL U1386 ( .A(n1548), .B(n1547), .Y(n1553) );
  NAND2XL U1387 ( .A(n1546), .B(n1549), .Y(n1556) );
  INVXL U1388 ( .A(n1550), .Y(n1546) );
  INVXL U1389 ( .A(n1554), .Y(n1561) );
  NAND2XL U1390 ( .A(n1539), .B(n1538), .Y(n1540) );
  NAND2BXL U1391 ( .AN(n1549), .B(n1550), .Y(n1538) );
  NAND2XL U1392 ( .A(n1550), .B(n1541), .Y(n1537) );
  NAND2XL U1393 ( .A(n1532), .B(n1531), .Y(n1539) );
  NAND2BXL U1394 ( .AN(n1527), .B(n1526), .Y(n1528) );
  NAND2XL U1395 ( .A(n1523), .B(n1522), .Y(n1529) );
  NAND2BXL U1396 ( .AN(n1519), .B(n1535), .Y(n1526) );
  NAND2XL U1397 ( .A(n1519), .B(n1520), .Y(n1524) );
  INVXL U1398 ( .A(n1505), .Y(n1507) );
  OAI211XL U1399 ( .A0(n1511), .A1(n1504), .B0(n1503), .C0(n1502), .Y(n1505)
         );
  INVXL U1400 ( .A(n1515), .Y(n1511) );
  NAND3XL U1401 ( .A(n1514), .B(n1517), .C(n1510), .Y(n1508) );
  NAND2XL U1402 ( .A(n1501), .B(n1500), .Y(n1510) );
  NOR2XL U1403 ( .A(n1501), .B(n1503), .Y(n1509) );
  NAND2XL U1404 ( .A(n1485), .B(n1483), .Y(n1494) );
  NOR2XL U1405 ( .A(n1489), .B(n1488), .Y(n1482) );
  INVXL U1406 ( .A(n1484), .Y(n1498) );
  NOR2BXL U1407 ( .AN(n173), .B(n1471), .Y(n1473) );
  NAND2XL U1408 ( .A(n1468), .B(n1469), .Y(n1477) );
  NAND2XL U1409 ( .A(n1471), .B(n173), .Y(n1469) );
  NAND4XL U1410 ( .A(n173), .B(n1472), .C(n1468), .D(n1467), .Y(n1464) );
  INVXL U1411 ( .A(n1476), .Y(n1468) );
  OAI2BB2XL U1412 ( .B0(next_work_cntr[19]), .B1(n1596), .A0N(
        next_work_cntr[19]), .A1N(n1596), .Y(n1470) );
  INVXL U1413 ( .A(next_work_cntr[6]), .Y(n1544) );
  NAND4XL U1414 ( .A(n1456), .B(n1455), .C(n1618), .D(n1621), .Y(n1612) );
  NOR4XL U1415 ( .A(n1719), .B(n1659), .C(n1640), .D(n1454), .Y(n1455) );
  NAND4XL U1416 ( .A(n1731), .B(n1738), .C(n1698), .D(n1678), .Y(n1454) );
  NAND2XL U1417 ( .A(n1383), .B(n898), .Y(n886) );
  INVXL U1418 ( .A(n1658), .Y(n1659) );
  INVXL U1419 ( .A(n1718), .Y(n1719) );
  NAND4XL U1420 ( .A(n1453), .B(n1652), .C(n1671), .D(n1633), .Y(n1613) );
  NOR2XL U1421 ( .A(n264), .B(n895), .Y(n896) );
  AOI211XL U1422 ( .A0(n1452), .A1(n1451), .B0(n1707), .C0(n1450), .Y(n1453)
         );
  OAI211XL U1423 ( .A0(N1184), .A1(n1778), .B0(n1753), .C0(n1691), .Y(n1450)
         );
  INVXL U1424 ( .A(n1747), .Y(n1753) );
  INVXL U1425 ( .A(n898), .Y(n1457) );
  NAND2XL U1426 ( .A(n360), .B(n606), .Y(n406) );
  NAND2XL U1427 ( .A(n360), .B(n591), .Y(n408) );
  NAND2XL U1428 ( .A(write_addr[6]), .B(n266), .Y(n409) );
  NAND2XL U1429 ( .A(n360), .B(n583), .Y(n411) );
  NAND2XL U1430 ( .A(n360), .B(n574), .Y(n413) );
  NAND2XL U1431 ( .A(n360), .B(n572), .Y(n414) );
  OAI211X1 U1432 ( .A0(n26), .A1(n1437), .B0(n1435), .C0(n1436), .Y(n2245) );
  AOI211XL U1433 ( .A0(n2225), .A1(n2235), .B0(n1434), .C0(n1940), .Y(n1437)
         );
  NAND2BXL U1434 ( .AN(n1411), .B(n1410), .Y(n1412) );
  OAI211XL U1435 ( .A0(n1423), .A1(n1409), .B0(n1408), .C0(n1419), .Y(n1410)
         );
  INVXL U1436 ( .A(n1419), .Y(n1425) );
  INVXL U1437 ( .A(n1392), .Y(n1390) );
  NAND2XL U1438 ( .A(n1385), .B(n1384), .Y(n1391) );
  NAND3XL U1439 ( .A(n1382), .B(n1388), .C(n1381), .Y(n1380) );
  NAND2XL U1440 ( .A(n1387), .B(n1386), .Y(n1382) );
  OAI211XL U1441 ( .A0(n1366), .A1(n1365), .B0(n1368), .C0(n1369), .Y(n1367)
         );
  NOR3XL U1442 ( .A(n1375), .B(n1377), .C(n175), .Y(n1372) );
  NOR2XL U1443 ( .A(n175), .B(n1376), .Y(n1373) );
  NAND2XL U1444 ( .A(n1364), .B(n1363), .Y(n1376) );
  INVXL U1445 ( .A(n1358), .Y(n1359) );
  NAND2BXL U1446 ( .AN(n1357), .B(n1369), .Y(n1362) );
  INVXL U1447 ( .A(n1355), .Y(n1365) );
  INVXL U1448 ( .A(n1352), .Y(n1354) );
  INVXL U1449 ( .A(n1843), .Y(n1847) );
  INVXL U1450 ( .A(n1846), .Y(n1863) );
  NAND2XL U1451 ( .A(n1352), .B(n1353), .Y(n1358) );
  INVXL U1452 ( .A(n1351), .Y(n1346) );
  OAI211XL U1453 ( .A0(n1351), .A1(n1352), .B0(n1347), .C0(n1341), .Y(n1345)
         );
  NAND2XL U1454 ( .A(n1340), .B(n1339), .Y(n1347) );
  INVXL U1455 ( .A(n1336), .Y(n1338) );
  NOR2XL U1456 ( .A(n1342), .B(n1341), .Y(n1332) );
  INVXL U1457 ( .A(n1328), .Y(n1329) );
  OAI211XL U1458 ( .A0(n1337), .A1(n1333), .B0(n1327), .C0(n1326), .Y(n1328)
         );
  INVXL U1459 ( .A(n1325), .Y(n1327) );
  NAND2XL U1460 ( .A(n1323), .B(n1322), .Y(n1331) );
  NAND2XL U1461 ( .A(n1318), .B(n1317), .Y(n1326) );
  NOR2XL U1462 ( .A(n1313), .B(n1318), .Y(n1315) );
  AOI32XL U1463 ( .A0(n1314), .A1(n1324), .A2(n1312), .B0(n1311), .B1(n1324), 
        .Y(n1316) );
  NAND2XL U1464 ( .A(n1310), .B(n1322), .Y(n1319) );
  NAND2XL U1465 ( .A(n1309), .B(n1308), .Y(n1322) );
  NAND2XL U1466 ( .A(n1298), .B(n1297), .Y(n1303) );
  NAND2XL U1467 ( .A(n1299), .B(n1300), .Y(n1312) );
  NAND4XL U1468 ( .A(n1293), .B(n1292), .C(n1298), .D(n1295), .Y(n1294) );
  NAND2XL U1469 ( .A(n1290), .B(n1293), .Y(n1297) );
  NOR2BXL U1470 ( .AN(n1293), .B(n1290), .Y(n1291) );
  INVXL U1471 ( .A(n1298), .Y(n1302) );
  INVXL U1472 ( .A(n1287), .Y(n1289) );
  NAND2XL U1473 ( .A(n622), .B(n621), .Y(n623) );
  INVXL U1474 ( .A(n620), .Y(n621) );
  NAND2XL U1475 ( .A(n1201), .B(n619), .Y(n624) );
  AND2XL U1476 ( .A(curr_photo_addr[19]), .B(n338), .Y(\C1/Z_19 ) );
  AOI211XL U1477 ( .A0(n613), .A1(n615), .B0(n612), .C0(n611), .Y(n614) );
  NOR2XL U1478 ( .A(n609), .B(n608), .Y(n612) );
  AOI211XL U1479 ( .A0(n150), .A1(n1974), .B0(n1973), .C0(n2211), .Y(n2048) );
  AOI211XL U1480 ( .A0(\next_write_addr_w[0] ), .A1(n1972), .B0(n150), .C0(
        n1971), .Y(n1973) );
  NOR2XL U1481 ( .A(n1972), .B(n1970), .Y(n1971) );
  NAND2XL U1482 ( .A(n2196), .B(n2045), .Y(n1974) );
  OAI211XL U1483 ( .A0(n2055), .A1(n2043), .B0(n659), .C0(n2057), .Y(n2044) );
  NOR2XL U1484 ( .A(n2127), .B(n149), .Y(n2046) );
  NAND2XL U1485 ( .A(read_cntr[1]), .B(n277), .Y(n424) );
  AOI211XL U1486 ( .A0(n355), .A1(n606), .B0(n605), .C0(n604), .Y(n607) );
  NOR2XL U1487 ( .A(n609), .B(n603), .Y(n605) );
  AOI211XL U1488 ( .A0(n613), .A1(n606), .B0(n601), .C0(n600), .Y(n602) );
  NOR2XL U1489 ( .A(n2233), .B(n608), .Y(n601) );
  OAI211XL U1490 ( .A0(write_addr[1]), .A1(write_addr[2]), .B0(n2090), .C0(
        n2066), .Y(n405) );
  AOI211XL U1491 ( .A0(n613), .A1(n598), .B0(n597), .C0(n596), .Y(n599) );
  NOR2XL U1492 ( .A(n593), .B(n608), .Y(n597) );
  INVXL U1493 ( .A(n2233), .Y(n598) );
  AND2XL U1494 ( .A(curr_photo_addr[5]), .B(n338), .Y(\C1/Z_5 ) );
  AOI211XL U1495 ( .A0(n355), .A1(n591), .B0(n590), .C0(n589), .Y(n592) );
  INVXL U1496 ( .A(n610), .Y(n595) );
  NOR2XL U1497 ( .A(n593), .B(n603), .Y(n590) );
  AND2XL U1498 ( .A(curr_photo_addr[6]), .B(n338), .Y(\C1/Z_6 ) );
  AOI211XL U1499 ( .A0(n613), .A1(n591), .B0(n587), .C0(n586), .Y(n588) );
  NOR2XL U1500 ( .A(n585), .B(n608), .Y(n587) );
  AOI211XL U1501 ( .A0(n355), .A1(n583), .B0(n582), .C0(n581), .Y(n584) );
  NOR2XL U1502 ( .A(n585), .B(n603), .Y(n582) );
  AND2XL U1503 ( .A(curr_photo_addr[8]), .B(n338), .Y(\C1/Z_8 ) );
  AOI211XL U1504 ( .A0(n613), .A1(n583), .B0(n578), .C0(n577), .Y(n580) );
  NOR2XL U1505 ( .A(n576), .B(n608), .Y(n578) );
  NOR2XL U1506 ( .A(n2110), .B(n2190), .Y(n2102) );
  AND2XL U1507 ( .A(curr_photo_addr[9]), .B(n338), .Y(\C1/Z_9 ) );
  AND2XL U1508 ( .A(curr_photo_addr[10]), .B(n338), .Y(\C1/Z_10 ) );
  AOI211XL U1509 ( .A0(n355), .A1(n572), .B0(n571), .C0(n570), .Y(n573) );
  NOR2XL U1510 ( .A(n576), .B(n603), .Y(n571) );
  AOI211XL U1511 ( .A0(n171), .A1(n2196), .B0(n2127), .C0(n149), .Y(n2103) );
  AOI211XL U1512 ( .A0(n613), .A1(n574), .B0(n568), .C0(n567), .Y(n569) );
  NOR2XL U1513 ( .A(n2229), .B(n608), .Y(n568) );
  XOR2XL U1514 ( .A(n2116), .B(n109), .Y(n412) );
  NOR2BXL U1515 ( .AN(n2115), .B(n2127), .Y(n2116) );
  AND2XL U1516 ( .A(curr_photo_addr[12]), .B(n338), .Y(\C1/Z_12 ) );
  AOI211XL U1517 ( .A0(n613), .A1(n572), .B0(n565), .C0(n564), .Y(n566) );
  NOR2XL U1518 ( .A(n563), .B(n608), .Y(n565) );
  AOI211XL U1519 ( .A0(n2129), .A1(n2128), .B0(n2174), .C0(n2211), .Y(n2130)
         );
  AOI211XL U1520 ( .A0(n613), .A1(n561), .B0(n560), .C0(n559), .Y(n562) );
  NOR2XL U1521 ( .A(n558), .B(n608), .Y(n560) );
  INVXL U1522 ( .A(n2229), .Y(n561) );
  INVXL U1523 ( .A(n2197), .Y(n2175) );
  AOI211XL U1524 ( .A0(n610), .A1(write_addr[12]), .B0(n556), .C0(n555), .Y(
        n557) );
  NOR2XL U1525 ( .A(n563), .B(n603), .Y(n556) );
  AOI211XL U1526 ( .A0(n2188), .A1(n2187), .B0(n2192), .C0(n2211), .Y(n2189)
         );
  AOI211XL U1527 ( .A0(n610), .A1(write_addr[13]), .B0(n552), .C0(n551), .Y(
        n553) );
  NOR2XL U1528 ( .A(n558), .B(n603), .Y(n552) );
  AOI211XL U1529 ( .A0(n2192), .A1(write_addr[13]), .B0(n2211), .C0(n416), .Y(
        n417) );
  NOR2XL U1530 ( .A(n2191), .B(n2192), .Y(n416) );
  NAND2XL U1531 ( .A(n109), .B(n2127), .Y(n2128) );
  OAI211XL U1532 ( .A0(n232), .A1(n2194), .B0(n659), .C0(n2193), .Y(n2195) );
  NAND2XL U1533 ( .A(n232), .B(n2194), .Y(n2186) );
  NAND3XL U1534 ( .A(n2184), .B(n2181), .C(n2183), .Y(n2182) );
  INVXL U1535 ( .A(n2180), .Y(n2183) );
  NOR2XL U1536 ( .A(n2123), .B(n2122), .Y(n2133) );
  AOI21XL U1537 ( .A0(n2121), .A1(n2120), .B0(\DP_OP_436J1_125_1438/n25 ), .Y(
        n2123) );
  NAND2BXL U1538 ( .AN(n170), .B(next_cr_x[6]), .Y(n333) );
  NAND2XL U1539 ( .A(next_cr_x[6]), .B(n170), .Y(n332) );
  NOR2XL U1540 ( .A(\DP_OP_436J1_125_1438/n26 ), .B(n2112), .Y(n2113) );
  NAND2BXL U1541 ( .AN(n2100), .B(n2099), .Y(n2108) );
  AND2XL U1542 ( .A(n2098), .B(\intadd_3/n1 ), .Y(n2097) );
  AOI22XL U1543 ( .A0(n2053), .A1(n2060), .B0(n2052), .B1(n2051), .Y(n2056) );
  NAND2XL U1544 ( .A(n2055), .B(n2043), .Y(n2057) );
  AOI21XL U1545 ( .A0(n2088), .A1(n2072), .B0(n2085), .Y(\intadd_3/B[0] ) );
  INVXL U1546 ( .A(n2068), .Y(\intadd_3/A[0] ) );
  INVXL U1547 ( .A(n2079), .Y(\intadd_3/B[1] ) );
  NAND2XL U1548 ( .A(n2064), .B(n2086), .Y(n2076) );
  INVXL U1549 ( .A(n2063), .Y(n2064) );
  NAND2XL U1550 ( .A(n2033), .B(n2032), .Y(n2038) );
  INVXL U1551 ( .A(n2035), .Y(n2028) );
  AOI22XL U1552 ( .A0(n177), .A1(n2022), .B0(n2026), .B1(n163), .Y(n2024) );
  AOI211XL U1553 ( .A0(n2078), .A1(n2021), .B0(n2020), .C0(n2019), .Y(n2022)
         );
  AOI21XL U1554 ( .A0(n2078), .A1(n2092), .B0(n2094), .Y(n2084) );
  AOI21XL U1555 ( .A0(n2083), .A1(n2082), .B0(n2106), .Y(n2093) );
  INVXL U1556 ( .A(n2013), .Y(n2016) );
  AND3XL U1557 ( .A(n2009), .B(n2008), .C(n2086), .Y(n2011) );
  NAND2XL U1558 ( .A(n2008), .B(n2086), .Y(n2007) );
  AOI21XL U1559 ( .A0(n2088), .A1(n2087), .B0(n2111), .Y(n2105) );
  INVXL U1560 ( .A(n1998), .Y(n2001) );
  NAND2XL U1561 ( .A(n2015), .B(n2010), .Y(n2014) );
  NAND3XL U1562 ( .A(n2012), .B(n2009), .C(n2008), .Y(n2010) );
  INVXL U1563 ( .A(n1993), .Y(n1994) );
  AND3XL U1564 ( .A(n1992), .B(n1991), .C(n2095), .Y(n1989) );
  INVXL U1565 ( .A(n1984), .Y(n1987) );
  NAND2XL U1566 ( .A(n2000), .B(n1988), .Y(n1999) );
  NAND3XL U1567 ( .A(n1992), .B(n1990), .C(n1991), .Y(n1988) );
  NAND2XL U1568 ( .A(n216), .B(n2107), .Y(n1993) );
  AND3XL U1569 ( .A(n1980), .B(n1979), .C(n2107), .Y(n1982) );
  INVXL U1570 ( .A(n909), .Y(n912) );
  NAND2XL U1571 ( .A(n1986), .B(n1981), .Y(n1985) );
  NAND3XL U1572 ( .A(n1983), .B(n1980), .C(n1979), .Y(n1981) );
  AND3XL U1573 ( .A(n903), .B(n902), .C(next_cr_x[5]), .Y(n900) );
  NOR2XL U1574 ( .A(n904), .B(next_cr_x[6]), .Y(n906) );
  AND2XL U1575 ( .A(next_cr_x[5]), .B(n170), .Y(n251) );
  AOI21XL U1576 ( .A0(n850), .A1(n2058), .B0(n2040), .Y(n853) );
  INVXL U1577 ( .A(n2053), .Y(n2062) );
  OAI211XL U1578 ( .A0(write_cntr[1]), .A1(write_cntr[0]), .B0(n845), .C0(n844), .Y(n846) );
  INVXL U1579 ( .A(n838), .Y(n842) );
  NAND4XL U1580 ( .A(write_cntr[1]), .B(n2040), .C(n849), .D(n2050), .Y(n855)
         );
  INVXL U1581 ( .A(n840), .Y(n843) );
  NAND2XL U1582 ( .A(n1443), .B(n2118), .Y(n835) );
  NAND2XL U1583 ( .A(n911), .B(n899), .Y(n910) );
  NAND3XL U1584 ( .A(n901), .B(n903), .C(n902), .Y(n899) );
  NAND2XL U1585 ( .A(next_cr_x[6]), .B(n904), .Y(n905) );
  INVXL U1586 ( .A(n1449), .Y(n728) );
  INVXL U1587 ( .A(n732), .Y(n709) );
  INVXL U1588 ( .A(n2119), .Y(n2118) );
  NOR2XL U1589 ( .A(n833), .B(n834), .Y(n831) );
  NOR2XL U1590 ( .A(n177), .B(n2172), .Y(n825) );
  NAND2XL U1591 ( .A(n824), .B(n823), .Y(n826) );
  NOR2XL U1592 ( .A(n2172), .B(n2180), .Y(n2173) );
  NAND2XL U1593 ( .A(n816), .B(n817), .Y(n815) );
  INVXL U1594 ( .A(n814), .Y(n817) );
  NOR2BXL U1595 ( .AN(n829), .B(n828), .Y(n818) );
  INVXL U1596 ( .A(n830), .Y(n828) );
  AOI21XL U1597 ( .A0(n813), .A1(n810), .B0(n812), .Y(n811) );
  NAND2XL U1598 ( .A(n2021), .B(n2170), .Y(n808) );
  NAND2XL U1599 ( .A(n824), .B(n1445), .Y(n819) );
  AOI221XL U1600 ( .A0(n270), .A1(n821), .B0(n149), .B1(n821), .C0(n807), .Y(
        n2023) );
  NOR2BXL U1601 ( .AN(n2171), .B(n2167), .Y(n2168) );
  NAND2XL U1602 ( .A(n2163), .B(n2162), .Y(n2165) );
  NAND2XL U1603 ( .A(n803), .B(n802), .Y(n814) );
  NAND2XL U1604 ( .A(n805), .B(n2163), .Y(n803) );
  NOR2XL U1605 ( .A(n2164), .B(n2017), .Y(n797) );
  NAND2XL U1606 ( .A(n796), .B(n800), .Y(n798) );
  INVXL U1607 ( .A(n722), .Y(n720) );
  NOR2XL U1608 ( .A(n2163), .B(n2162), .Y(n2160) );
  NOR2BXL U1609 ( .AN(n2166), .B(n2164), .Y(n2161) );
  NAND2XL U1610 ( .A(n2156), .B(n2155), .Y(n2158) );
  NAND3XL U1611 ( .A(n2156), .B(n2159), .C(n2155), .Y(n2154) );
  AND2XL U1612 ( .A(n2150), .B(n2152), .Y(n2151) );
  NAND2XL U1613 ( .A(n2150), .B(n2152), .Y(n2148) );
  NAND2XL U1614 ( .A(n2152), .B(n2153), .Y(n2149) );
  NAND2XL U1615 ( .A(n2144), .B(n2143), .Y(n2146) );
  NAND3XL U1616 ( .A(n2144), .B(n2147), .C(n2143), .Y(n2142) );
  NAND3XL U1617 ( .A(n2141), .B(n237), .C(n2140), .Y(n2139) );
  NAND2XL U1618 ( .A(n2140), .B(n2141), .Y(n2137) );
  NAND2XL U1619 ( .A(n793), .B(n794), .Y(n792) );
  INVXL U1620 ( .A(n791), .Y(n794) );
  NOR2BXL U1621 ( .AN(n805), .B(n804), .Y(n795) );
  INVXL U1622 ( .A(n806), .Y(n804) );
  AOI21XL U1623 ( .A0(n790), .A1(n787), .B0(n789), .Y(n788) );
  NAND2XL U1624 ( .A(n2002), .B(n796), .Y(n801) );
  NAND2XL U1625 ( .A(n782), .B(n784), .Y(n781) );
  INVXL U1626 ( .A(n780), .Y(n782) );
  NOR2XL U1627 ( .A(n793), .B(n791), .Y(n785) );
  NOR2XL U1628 ( .A(n783), .B(n216), .Y(n774) );
  NAND2XL U1629 ( .A(n784), .B(n780), .Y(n772) );
  NAND2XL U1630 ( .A(n1444), .B(n2143), .Y(n767) );
  NOR2XL U1631 ( .A(n770), .B(n771), .Y(n761) );
  INVXL U1632 ( .A(n760), .Y(n765) );
  NAND2XL U1633 ( .A(n753), .B(n754), .Y(n752) );
  INVXL U1634 ( .A(n751), .Y(n753) );
  NOR2XL U1635 ( .A(n904), .B(n2138), .Y(n749) );
  INVXL U1636 ( .A(n755), .Y(n764) );
  NAND2XL U1637 ( .A(n1444), .B(n768), .Y(n755) );
  INVXL U1638 ( .A(n242), .Y(n747) );
  NAND2XL U1639 ( .A(n908), .B(n2136), .Y(n739) );
  NAND2XL U1640 ( .A(n1446), .B(n750), .Y(n748) );
  NAND2BXL U1641 ( .AN(n746), .B(n242), .Y(n736) );
  INVXL U1642 ( .A(n731), .Y(n733) );
  NAND2XL U1643 ( .A(n254), .B(n702), .Y(n701) );
  NAND2XL U1644 ( .A(n716), .B(n715), .Y(n717) );
  NAND4XL U1645 ( .A(write_cntr[7]), .B(write_cntr[6]), .C(write_cntr[8]), .D(
        n724), .Y(n716) );
  NAND2XL U1646 ( .A(n220), .B(n727), .Y(n726) );
  NAND3XL U1647 ( .A(write_cntr[6]), .B(n724), .C(n845), .Y(n727) );
  INVXL U1648 ( .A(n837), .Y(n845) );
  NOR2XL U1649 ( .A(n837), .B(n723), .Y(n725) );
  INVXL U1650 ( .A(n724), .Y(n723) );
  NAND2XL U1651 ( .A(n253), .B(n722), .Y(n721) );
  NAND3XL U1652 ( .A(write_cntr[4]), .B(write_cntr[3]), .C(write_cntr[2]), .Y(
        n719) );
  NOR2XL U1653 ( .A(n245), .B(n714), .Y(n698) );
  NAND2XL U1654 ( .A(write_cntr[7]), .B(write_cntr[6]), .Y(n714) );
  AND2XL U1655 ( .A(curr_photo_addr[16]), .B(n338), .Y(\C1/Z_16 ) );
  AOI211XL U1656 ( .A0(write_addr[14]), .A1(n610), .B0(n548), .C0(n547), .Y(
        n549) );
  NOR2XL U1657 ( .A(n603), .B(n554), .Y(n548) );
  AND2XL U1658 ( .A(curr_photo_addr[17]), .B(n338), .Y(\C1/Z_17 ) );
  AOI211XL U1659 ( .A0(write_addr[15]), .A1(n610), .B0(n545), .C0(n544), .Y(
        n546) );
  NOR2XL U1660 ( .A(n603), .B(n550), .Y(n545) );
  XNOR2XL U1661 ( .A(write_addr[15]), .B(n2202), .Y(n418) );
  NAND2XL U1662 ( .A(write_addr[14]), .B(n2201), .Y(n2202) );
  AND2XL U1663 ( .A(curr_photo_addr[18]), .B(n338), .Y(\C1/Z_18 ) );
  AOI211XL U1664 ( .A0(write_addr[16]), .A1(n610), .B0(n542), .C0(n541), .Y(
        n543) );
  INVXL U1665 ( .A(n2208), .Y(n2209) );
  NOR2XL U1666 ( .A(n2231), .B(n603), .Y(n542) );
  NAND2XL U1667 ( .A(write_addr[16]), .B(n2206), .Y(n2208) );
  OAI21X1 U1668 ( .A0(n661), .A1(n693), .B0(n691), .Y(next_state[2]) );
  OA21X4 U1669 ( .A0(n696), .A1(n26), .B0(n697), .Y(n220) );
  AOI22X1 U1670 ( .A0(n26), .A1(n689), .B0(n234), .B1(n691), .Y(n697) );
  OAI21X1 U1671 ( .A0(n26), .A1(n2218), .B0(n688), .Y(n691) );
  INVXL U1672 ( .A(n687), .Y(n688) );
  NAND2XL U1673 ( .A(n678), .B(n670), .Y(n690) );
  OAI211XL U1674 ( .A0(n669), .A1(n674), .B0(n641), .C0(n107), .Y(n670) );
  AOI211XL U1675 ( .A0(n667), .A1(n666), .B0(n672), .C0(n250), .Y(n669) );
  INVXL U1676 ( .A(n647), .Y(n672) );
  INVXL U1677 ( .A(n1614), .Y(n683) );
  INVXL U1678 ( .A(n694), .Y(n661) );
  NAND4XL U1679 ( .A(n678), .B(n677), .C(n676), .D(n675), .Y(n679) );
  NOR4XL U1680 ( .A(n647), .B(n646), .C(n649), .D(n674), .Y(n675) );
  NOR4XL U1681 ( .A(n653), .B(n650), .C(n655), .D(n654), .Y(n676) );
  AOI21X1 U1682 ( .A0(n241), .A1(n362), .B0(n652), .Y(n653) );
  NOR2XL U1683 ( .A(n651), .B(next_glb_cntr[6]), .Y(n677) );
  NAND3XL U1684 ( .A(n652), .B(n665), .C(n246), .Y(n363) );
  NAND2XL U1685 ( .A(global_cntr[17]), .B(n372), .Y(n373) );
  XNOR2XL U1686 ( .A(n372), .B(n107), .Y(n371) );
  NAND2BXL U1687 ( .AN(n665), .B(n652), .Y(n671) );
  NOR2X2 U1688 ( .A(n362), .B(n241), .Y(n652) );
  NAND2X1 U1689 ( .A(n361), .B(global_cntr[4]), .Y(n362) );
  NAND3XL U1690 ( .A(global_cntr[17]), .B(global_cntr[18]), .C(global_cntr[16]), .Y(n662) );
  NOR3XL U1691 ( .A(n2197), .B(n171), .C(n2196), .Y(n2198) );
  AOI211XL U1692 ( .A0(n1967), .A1(n2213), .B0(n1966), .C0(n2101), .Y(n2049)
         );
  AOI211XL U1693 ( .A0(write_addr[4]), .A1(n2075), .B0(n2091), .C0(n630), .Y(
        n1966) );
  NOR4XL U1694 ( .A(n2210), .B(n2214), .C(n2207), .D(n1961), .Y(n1967) );
  AOI21XL U1695 ( .A0(n2197), .A1(n2188), .B0(n2205), .Y(n1961) );
  AND2XL U1696 ( .A(n1956), .B(write_addr[17]), .Y(n1962) );
  NAND3XL U1697 ( .A(write_addr[15]), .B(write_addr[14]), .C(n2191), .Y(n2205)
         );
  INVXL U1698 ( .A(n2125), .Y(n1958) );
  NAND2XL U1699 ( .A(n2126), .B(write_addr[10]), .Y(n2125) );
  NAND2XL U1700 ( .A(n1965), .B(write_addr[7]), .Y(n1964) );
  AND2XL U1701 ( .A(n1963), .B(write_addr[6]), .Y(n1965) );
  NAND2XL U1702 ( .A(n2227), .B(n2226), .Y(n2228) );
  NAND2XL U1703 ( .A(n2223), .B(n2236), .Y(n2234) );
  NOR2XL U1704 ( .A(read_cntr[0]), .B(read_cntr[1]), .Y(n2227) );
  NAND2XL U1705 ( .A(n619), .B(n632), .Y(n399) );
  NAND2BXL U1706 ( .AN(n2236), .B(n1911), .Y(n619) );
  INVXL U1707 ( .A(n1201), .Y(n400) );
  NOR2XL U1708 ( .A(n1200), .B(n1199), .Y(n1198) );
  NAND2XL U1709 ( .A(n1452), .B(n1197), .Y(n1191) );
  NAND2XL U1710 ( .A(n1783), .B(n1190), .Y(n1452) );
  NOR2XL U1711 ( .A(n1192), .B(n2235), .Y(n1193) );
  INVXL U1712 ( .A(n1186), .Y(n1196) );
  NAND3XL U1713 ( .A(n1183), .B(n1180), .C(n1182), .Y(n1181) );
  NOR2BXL U1714 ( .AN(n1188), .B(n1756), .Y(n1185) );
  NAND3XL U1715 ( .A(n1170), .B(n1169), .C(n1165), .Y(n1168) );
  INVXL U1716 ( .A(n1173), .Y(n1167) );
  INVXL U1717 ( .A(n1157), .Y(n1158) );
  INVXL U1718 ( .A(n1166), .Y(n1175) );
  NOR2XL U1719 ( .A(work_cntr[4]), .B(n1171), .Y(n1153) );
  INVXL U1720 ( .A(n1163), .Y(n1164) );
  NAND3XL U1721 ( .A(n1157), .B(n1151), .C(n1154), .Y(n1165) );
  NAND3XL U1722 ( .A(n1156), .B(n1155), .C(n1150), .Y(n1154) );
  INVXL U1723 ( .A(n1149), .Y(n1155) );
  AOI21XL U1724 ( .A0(n265), .A1(n1149), .B0(n1144), .Y(n1145) );
  INVXL U1725 ( .A(n1151), .Y(n1160) );
  NOR2BXL U1726 ( .AN(n1140), .B(work_cntr[7]), .Y(n1139) );
  NAND3XL U1727 ( .A(n1144), .B(n204), .C(n1141), .Y(n1150) );
  NAND3XL U1728 ( .A(n1143), .B(n1142), .C(n1137), .Y(n1141) );
  INVXL U1729 ( .A(n1143), .Y(n1133) );
  INVXL U1730 ( .A(n1135), .Y(n1142) );
  INVXL U1731 ( .A(n1130), .Y(n1132) );
  NAND3XL U1732 ( .A(n1123), .B(n1129), .C(n1125), .Y(n1137) );
  NAND3XL U1733 ( .A(n1127), .B(n1126), .C(n1122), .Y(n1125) );
  INVXL U1734 ( .A(n1121), .Y(n1127) );
  INVXL U1735 ( .A(n1128), .Y(n1123) );
  INVXL U1736 ( .A(n1114), .Y(n1115) );
  INVXL U1737 ( .A(n1119), .Y(n1120) );
  INVXL U1738 ( .A(n1113), .Y(n1106) );
  NAND2XL U1739 ( .A(n1097), .B(n1096), .Y(n1101) );
  INVXL U1740 ( .A(n1093), .Y(n1095) );
  NOR2XL U1741 ( .A(work_cntr[12]), .B(n1107), .Y(n1091) );
  NOR2XL U1742 ( .A(n1109), .B(n1103), .Y(n1104) );
  INVXL U1743 ( .A(n211), .Y(n1086) );
  NAND2XL U1744 ( .A(n1082), .B(n1798), .Y(n1093) );
  NAND2XL U1745 ( .A(n1083), .B(n1094), .Y(n1088) );
  NAND2XL U1746 ( .A(n1078), .B(n1077), .Y(n1079) );
  NAND2XL U1747 ( .A(work_cntr[17]), .B(n1084), .Y(n1081) );
  NAND2BXL U1748 ( .AN(n1078), .B(work_cntr[18]), .Y(n1076) );
  INVXL U1749 ( .A(n1089), .Y(n1099) );
  INVXL U1750 ( .A(n1074), .Y(n1075) );
  INVXL U1751 ( .A(n1414), .Y(n1451) );
  NAND3X1 U1752 ( .A(en_so), .B(n26), .C(n1933), .Y(n620) );
  NAND2BX4 U1753 ( .AN(n694), .B(n687), .Y(en_so) );
  NAND2XL U1754 ( .A(n1072), .B(n1073), .Y(n398) );
  AOI22XL U1755 ( .A0(n1068), .A1(n1067), .B0(n1066), .B1(n1065), .Y(n1071) );
  NAND2BXL U1756 ( .AN(n1065), .B(n1063), .Y(n1062) );
  MXI2XL U1757 ( .A(n1066), .B(n1065), .S0(n1063), .Y(n1068) );
  NAND2XL U1758 ( .A(n1073), .B(n1069), .Y(n1070) );
  NOR2XL U1759 ( .A(n1066), .B(n1063), .Y(n1061) );
  INVXL U1760 ( .A(n1056), .Y(n1060) );
  INVXL U1761 ( .A(n1057), .Y(n1053) );
  NOR2XL U1762 ( .A(N1183), .B(n1056), .Y(n1052) );
  NAND2XL U1763 ( .A(n1057), .B(n1051), .Y(n1055) );
  INVXL U1764 ( .A(n1046), .Y(n1044) );
  INVXL U1765 ( .A(n1043), .Y(n1048) );
  NAND2XL U1766 ( .A(n1042), .B(n1046), .Y(n1050) );
  NAND2XL U1767 ( .A(n1041), .B(n1040), .Y(n1046) );
  INVXL U1768 ( .A(n1034), .Y(n1038) );
  NOR2XL U1769 ( .A(N1184), .B(n1043), .Y(n1039) );
  NOR2XL U1770 ( .A(work_cntr[4]), .B(n1034), .Y(n1033) );
  NAND2XL U1771 ( .A(n160), .B(n1035), .Y(n1040) );
  NAND2XL U1772 ( .A(n1029), .B(n1031), .Y(n1035) );
  NAND2BXL U1773 ( .AN(n1028), .B(n1027), .Y(n1031) );
  NAND2XL U1774 ( .A(n1024), .B(n1023), .Y(n1027) );
  NAND2XL U1775 ( .A(n1022), .B(n1028), .Y(n1029) );
  NAND2XL U1776 ( .A(n1020), .B(n1018), .Y(n1019) );
  NAND2XL U1777 ( .A(n1026), .B(n229), .Y(n1022) );
  NOR2XL U1778 ( .A(work_cntr[6]), .B(n1020), .Y(n1017) );
  NAND2XL U1779 ( .A(n1016), .B(n1021), .Y(n1023) );
  NAND2XL U1780 ( .A(n1012), .B(n1011), .Y(n1015) );
  NAND2XL U1781 ( .A(n1008), .B(n1007), .Y(n1011) );
  NOR2XL U1782 ( .A(work_cntr[7]), .B(n1005), .Y(n1006) );
  INVXL U1783 ( .A(n1005), .Y(n1010) );
  NAND2XL U1784 ( .A(n1000), .B(n999), .Y(n1008) );
  NAND2XL U1785 ( .A(n1004), .B(n262), .Y(n1000) );
  NAND2BXL U1786 ( .AN(n999), .B(n1001), .Y(n1007) );
  NAND2XL U1787 ( .A(n995), .B(n994), .Y(n998) );
  NAND2XL U1788 ( .A(n993), .B(n997), .Y(n992) );
  INVXL U1789 ( .A(n994), .Y(n991) );
  INVXL U1790 ( .A(n985), .Y(n989) );
  NOR2XL U1791 ( .A(work_cntr[9]), .B(n993), .Y(n990) );
  INVXL U1792 ( .A(n986), .Y(n982) );
  NAND2XL U1793 ( .A(n981), .B(n986), .Y(n984) );
  NAND2XL U1794 ( .A(n980), .B(n979), .Y(n986) );
  NOR2XL U1795 ( .A(work_cntr[10]), .B(n985), .Y(n978) );
  NAND2BXL U1796 ( .AN(n976), .B(n975), .Y(n979) );
  NAND2XL U1797 ( .A(n976), .B(n970), .Y(n980) );
  NAND2XL U1798 ( .A(n974), .B(n267), .Y(n970) );
  NAND2XL U1799 ( .A(n968), .B(n966), .Y(n967) );
  INVXL U1800 ( .A(n969), .Y(n965) );
  NOR2XL U1801 ( .A(work_cntr[12]), .B(n968), .Y(n963) );
  NAND2XL U1802 ( .A(n964), .B(n969), .Y(n971) );
  NAND2XL U1803 ( .A(n959), .B(n958), .Y(n962) );
  INVXL U1804 ( .A(n958), .Y(n955) );
  NAND2XL U1805 ( .A(n957), .B(n268), .Y(n952) );
  NAND3XL U1806 ( .A(n946), .B(n943), .C(n264), .Y(n944) );
  NOR2XL U1807 ( .A(work_cntr[15]), .B(n947), .Y(n945) );
  NAND2XL U1808 ( .A(n946), .B(n264), .Y(n940) );
  INVXL U1809 ( .A(n936), .Y(n937) );
  NOR2XL U1810 ( .A(work_cntr[17]), .B(n1619), .Y(n938) );
  INVXL U1811 ( .A(n1792), .Y(n1619) );
  INVXL U1812 ( .A(n1077), .Y(n1626) );
  NAND2XL U1813 ( .A(n934), .B(n260), .Y(n936) );
  INVXL U1814 ( .A(n1286), .Y(n935) );
  OAI211XL U1815 ( .A0(work_cntr[16]), .A1(n236), .B0(work_cntr[17]), .C0(n259), .Y(n933) );
  NOR4XL U1816 ( .A(N76), .B(n1433), .C(n1432), .D(n1431), .Y(n1434) );
  MXI2XL U1817 ( .A(n1951), .B(n1942), .S0(N684), .Y(n316) );
  AND3XL U1818 ( .A(N684), .B(N685), .C(n1947), .Y(n631) );
  NOR4XL U1819 ( .A(n662), .B(n233), .C(n243), .D(n926), .Y(n663) );
  OAI22XL U1820 ( .A0(n622), .A1(n620), .B0(n400), .B1(n399), .Y(
        \RSOP_434/C2/CONTROL1 ) );
  NOR2XL U1821 ( .A(N76), .B(n1064), .Y(n1072) );
  NAND2XL U1822 ( .A(N76), .B(n1064), .Y(n1067) );
  NOR3BX1 U1823 ( .AN(n930), .B(global_cntr[19]), .C(n929), .Y(n1282) );
  NAND4XL U1824 ( .A(n928), .B(n927), .C(n247), .D(n225), .Y(n929) );
  NOR4XL U1825 ( .A(global_cntr[3]), .B(global_cntr[4]), .C(n926), .D(n925), 
        .Y(n927) );
  OAI22XL U1826 ( .A0(n2222), .A1(n423), .B0(n2221), .B1(n325), .Y(
        next_photo[1]) );
  OAI21XL U1827 ( .A0(cr_read_cntr[3]), .A1(n535), .B0(n536), .Y(N29) );
  AO22X1 U1828 ( .A0(write_addr[18]), .A1(n266), .B0(n540), .B1(n420), .Y(n289) );
  AOI211XL U1829 ( .A0(n1427), .A1(n257), .B0(n228), .C0(n1426), .Y(n1428) );
  NAND2BX1 U1830 ( .AN(n2242), .B(n2241), .Y(so_mux_sel[1]) );
  AO21X1 U1831 ( .A0(n632), .A1(n2240), .B0(n2242), .Y(so_mux_sel[0]) );
  OAI31XL U1832 ( .A0(n2237), .A1(n2236), .A2(n2235), .B0(n2234), .Y(n2240) );
  OAI22XL U1833 ( .A0(n360), .A1(n276), .B0(n539), .B1(im_wen_n), .Y(n288) );
  OAI22XL U1834 ( .A0(n360), .A1(n2230), .B0(n2231), .B1(im_wen_n), .Y(n291)
         );
  OAI22XL U1835 ( .A0(n360), .A1(n274), .B0(n554), .B1(im_wen_n), .Y(n293) );
  OAI22XL U1836 ( .A0(n360), .A1(n2203), .B0(im_wen_n), .B1(n550), .Y(n292) );
  OAI22XL U1837 ( .A0(n360), .A1(n318), .B0(n2232), .B1(im_wen_n), .Y(n290) );
  OAI22XL U1838 ( .A0(n147), .A1(n729), .B0(n360), .B1(n324), .Y(n340) );
  OAI22XL U1839 ( .A0(n147), .A1(n1445), .B0(n360), .B1(n270), .Y(n348) );
  OAI22XL U1840 ( .A0(n147), .A1(n1978), .B0(n360), .B1(n256), .Y(n345) );
  OAI22XL U1841 ( .A0(n147), .A1(n2002), .B0(n360), .B1(n253), .Y(n347) );
  OAI22XL U1842 ( .A0(n147), .A1(n1444), .B0(n360), .B1(n245), .Y(n351) );
  OAI22XL U1843 ( .A0(n230), .A1(n360), .B0(n1446), .B1(im_wen_n), .Y(n344) );
  OAI22XL U1844 ( .A0(n254), .A1(n360), .B0(n1449), .B1(im_wen_n), .Y(n339) );
  OAI22XL U1845 ( .A0(n248), .A1(n360), .B0(n1447), .B1(im_wen_n), .Y(n342) );
  OAI22XL U1846 ( .A0(n147), .A1(n908), .B0(n360), .B1(n113), .Y(n343) );
  OAI22XL U1847 ( .A0(n285), .A1(n360), .B0(n2021), .B1(im_wen_n), .Y(n352) );
  OAI2BB2XL U1848 ( .B0(n360), .B1(n271), .A0N(n360), .A1N(n1442), .Y(n354) );
  OAI22XL U1849 ( .A0(n2243), .A1(n326), .B0(n425), .B1(n2244), .Y(n335) );
  AOI21XL U1850 ( .A0(N684), .A1(n1947), .B0(N685), .Y(n401) );
  OAI21XL U1851 ( .A0(n1941), .A1(n224), .B0(n402), .Y(n314) );
  OAI21XL U1852 ( .A0(n360), .A1(n330), .B0(n422), .Y(n307) );
  OAI21XL U1853 ( .A0(n609), .A1(n266), .B0(n404), .Y(n306) );
  NOR4XL U1854 ( .A(n323), .B(n231), .C(n240), .D(n224), .Y(n1943) );
  OAI21XL U1855 ( .A0(n360), .A1(n329), .B0(n406), .Y(n305) );
  OAI21XL U1856 ( .A0(n360), .A1(n239), .B0(n408), .Y(n302) );
  OAI21XL U1857 ( .A0(n585), .A1(n266), .B0(n409), .Y(n301) );
  OAI21XL U1858 ( .A0(n360), .A1(n328), .B0(n411), .Y(n300) );
  OAI21XL U1859 ( .A0(n360), .A1(n273), .B0(n413), .Y(n298) );
  OAI21XL U1860 ( .A0(n360), .A1(n327), .B0(n414), .Y(n297) );
  OAI21XL U1861 ( .A0(n563), .A1(n147), .B0(n415), .Y(n295) );
  NOR2X1 U1862 ( .A(n637), .B(n338), .Y(n1436) );
  CLKBUFX3 U1863 ( .A(n625), .Y(n356) );
  AOI2BB1X1 U1864 ( .A0N(n2193), .A1N(n2190), .B0(n2189), .Y(n563) );
  OAI31XL U1865 ( .A0(write_cntr[9]), .A1(write_cntr[10]), .A2(n698), .B0(
        write_cntr[11]), .Y(n699) );
  NOR3XL U1866 ( .A(write_cntr[14]), .B(write_cntr[13]), .C(write_cntr[12]), 
        .Y(n700) );
  CLKINVX1 U1867 ( .A(n695), .Y(n2219) );
  CLKINVX1 U1868 ( .A(n632), .Y(n2238) );
  CLKINVX1 U1869 ( .A(n2211), .Y(n660) );
  NOR2X1 U1870 ( .A(next_state[2]), .B(next_state[1]), .Y(n695) );
  AO22X1 U1871 ( .A0(n694), .A1(n693), .B0(n48), .B1(n692), .Y(next_state[1])
         );
  NAND2XL U1872 ( .A(n252), .B(n690), .Y(n693) );
  OAI21XL U1873 ( .A0(n924), .A1(n683), .B0(n337), .Y(n684) );
  NOR2X1 U1874 ( .A(n248), .B(n682), .Y(n1936) );
  NAND4XL U1875 ( .A(write_cntr[13]), .B(write_cntr[14]), .C(write_cntr[12]), 
        .D(n681), .Y(n682) );
  AOI21XL U1876 ( .A0(global_cntr[6]), .A1(n652), .B0(global_cntr[7]), .Y(n364) );
  XNOR2XL U1877 ( .A(n664), .B(global_cntr[19]), .Y(n374) );
  NOR2X1 U1878 ( .A(n244), .B(n367), .Y(n368) );
  NAND4XL U1879 ( .A(n928), .B(n930), .C(global_cntr[19]), .D(n663), .Y(n665)
         );
  OR2X4 U1880 ( .A(\DP_OP_438J1_134_2124/I5 ), .B(si_sel), .Y(n626) );
  OR2X4 U1881 ( .A(n338), .B(n48), .Y(\DP_OP_438J1_134_2124/I5 ) );
  NAND2X1 U1882 ( .A(n1413), .B(n1172), .Y(n2236) );
  CLKINVX1 U1883 ( .A(n1429), .Y(n1413) );
  NOR2X1 U1884 ( .A(n2190), .B(n1940), .Y(n1938) );
  NAND2X1 U1885 ( .A(n690), .B(n687), .Y(n686) );
  AOI21X1 U1886 ( .A0(n244), .A1(n367), .B0(n368), .Y(n645) );
  NOR2X1 U1887 ( .A(n225), .B(n668), .Y(n372) );
  NOR2X1 U1888 ( .A(n243), .B(n369), .Y(n370) );
  CLKINVX1 U1889 ( .A(n932), .Y(n377) );
  NOR2X1 U1890 ( .A(work_cntr[19]), .B(n1286), .Y(n1793) );
  AOI2BB1X1 U1891 ( .A0N(global_cntr[1]), .A1N(global_cntr[0]), .B0(n657), .Y(
        next_glb_cntr[1]) );
  OAI22XL U1892 ( .A0(n487), .A1(n486), .B0(n485), .B1(n484), .Y(n488) );
  OAI21XL U1893 ( .A0(n882), .A1(n460), .B0(n459), .Y(n461) );
  AOI2BB2X1 U1894 ( .B0(n517), .B1(n465), .A0N(n532), .A1N(n451), .Y(n494) );
  AOI2BB2X1 U1895 ( .B0(n529), .B1(n507), .A0N(n879), .A1N(n527), .Y(n508) );
  OAI21XL U1896 ( .A0(n512), .A1(n506), .B0(n505), .Y(n507) );
  OAI21XL U1897 ( .A0(curr_time[9]), .A1(n512), .B0(n504), .Y(n505) );
  OR2X1 U1898 ( .A(curr_time[9]), .B(n504), .Y(n506) );
  OAI21XL U1899 ( .A0(n502), .A1(n501), .B0(n500), .Y(n503) );
  AOI2BB2X1 U1900 ( .B0(n518), .B1(n499), .A0N(n531), .A1N(n498), .Y(n510) );
  OAI21XL U1901 ( .A0(n497), .A1(n496), .B0(n495), .Y(n499) );
  OAI21XL U1902 ( .A0(n445), .A1(n441), .B0(curr_time[18]), .Y(n442) );
  OAI21XL U1903 ( .A0(n881), .A1(n658), .B0(n455), .Y(n457) );
  OAI2BB1X1 U1904 ( .A0N(n396), .A1N(n395), .B0(n394), .Y(n460) );
  AOI2BB2X1 U1905 ( .B0(n393), .B1(n392), .A0N(n877), .A1N(n878), .Y(n397) );
  AOI2BB2X1 U1906 ( .B0(n862), .B1(n436), .A0N(n435), .A1N(n863), .Y(n439) );
  OAI2BB1X1 U1907 ( .A0N(n435), .A1N(n434), .B0(n433), .Y(n440) );
  OR2X1 U1908 ( .A(n432), .B(n431), .Y(n443) );
  OAI2BB1X1 U1909 ( .A0N(n476), .A1N(n475), .B0(n474), .Y(n485) );
  OAI2BB1X1 U1910 ( .A0N(n473), .A1N(n472), .B0(n471), .Y(n479) );
  OR2X1 U1911 ( .A(n169), .B(n1440), .Y(n532) );
  NAND3BX1 U1912 ( .AN(n1439), .B(n1277), .C(n426), .Y(n452) );
  OA21XL U1913 ( .A0(n538), .A1(n537), .B0(n536), .Y(N28) );
  AND2XL U1914 ( .A(n1427), .B(n257), .Y(n1416) );
  OA21XL U1915 ( .A0(cr_read_cntr[3]), .A1(n403), .B0(n1945), .Y(n313) );
  OAI211XL U1916 ( .A0(n1924), .A1(n227), .B0(n1925), .C0(n257), .Y(n1923) );
  NOR2XL U1917 ( .A(N1182), .B(N1183), .Y(n1912) );
  NAND2X1 U1918 ( .A(write_addr[12]), .B(n147), .Y(n415) );
  CLKINVX1 U1919 ( .A(en_so), .Y(n637) );
  OAI22XL U1920 ( .A0(n618), .A1(n614), .B0(n334), .B1(n249), .Y(\C2/Z_1 ) );
  AO22X1 U1921 ( .A0(n610), .A1(\next_write_addr_w[0] ), .B0(n616), .B1(
        write_addr[1]), .Y(n611) );
  AO22X1 U1922 ( .A0(curr_photo_addr[1]), .A1(n338), .B0(n48), .B1(
        curr_photo[0]), .Y(n627) );
  OR2X1 U1923 ( .A(n2047), .B(n2048), .Y(n615) );
  AO22X1 U1924 ( .A0(curr_photo_addr[2]), .A1(n338), .B0(n48), .B1(
        curr_photo[1]), .Y(n628) );
  OAI22XL U1925 ( .A0(n618), .A1(n607), .B0(n334), .B1(n226), .Y(\C2/Z_2 ) );
  AO22X1 U1926 ( .A0(n610), .A1(write_addr[1]), .B0(n616), .B1(write_addr[2]), 
        .Y(n604) );
  OA22X1 U1927 ( .A0(n2190), .A1(n2054), .B0(write_addr[1]), .B1(n410), .Y(
        n609) );
  AO21X1 U1928 ( .A0(curr_photo_addr[3]), .A1(n338), .B0(si_sel), .Y(n629) );
  OAI22XL U1929 ( .A0(n618), .A1(n602), .B0(n334), .B1(n280), .Y(\C2/Z_3 ) );
  AO22X1 U1930 ( .A0(n610), .A1(write_addr[2]), .B0(n616), .B1(write_addr[3]), 
        .Y(n600) );
  AO21X1 U1931 ( .A0(curr_photo_addr[4]), .A1(n338), .B0(si_sel), .Y(\C1/Z_4 )
         );
  OAI22XL U1932 ( .A0(n618), .A1(n599), .B0(n334), .B1(n282), .Y(\C2/Z_4 ) );
  OAI22XL U1933 ( .A0(n595), .A1(n238), .B0(n594), .B1(n281), .Y(n596) );
  OAI22XL U1934 ( .A0(n618), .A1(n592), .B0(n334), .B1(n241), .Y(\C2/Z_5 ) );
  OAI22XL U1935 ( .A0(n595), .A1(n281), .B0(n594), .B1(n239), .Y(n589) );
  AOI2BB2X1 U1936 ( .B0(\intadd_3/SUM[1] ), .B1(n659), .A0N(n407), .A1N(n410), 
        .Y(n593) );
  OAI21XL U1937 ( .A0(n2080), .A1(write_addr[4]), .B0(n2081), .Y(n407) );
  OAI22XL U1938 ( .A0(n618), .A1(n588), .B0(n334), .B1(n246), .Y(\C2/Z_6 ) );
  AO22X1 U1939 ( .A0(n610), .A1(write_addr[5]), .B0(n616), .B1(write_addr[6]), 
        .Y(n586) );
  AO22X1 U1940 ( .A0(\intadd_3/SUM[2] ), .A1(n659), .B0(n630), .B1(n2090), .Y(
        n591) );
  AO21X1 U1941 ( .A0(curr_photo_addr[7]), .A1(n338), .B0(si_sel), .Y(\C1/Z_7 )
         );
  OAI22XL U1942 ( .A0(n618), .A1(n584), .B0(n334), .B1(n283), .Y(\C2/Z_7 ) );
  AO22X1 U1943 ( .A0(n610), .A1(write_addr[6]), .B0(n616), .B1(write_addr[7]), 
        .Y(n581) );
  AOI2BB2X1 U1944 ( .B0(n2090), .B1(n2091), .A0N(n2097), .A1N(n2089), .Y(n585)
         );
  OAI22XL U1945 ( .A0(n618), .A1(n580), .B0(n334), .B1(n579), .Y(\C2/Z_8 ) );
  AO22X1 U1946 ( .A0(n610), .A1(write_addr[7]), .B0(n616), .B1(n112), .Y(n577)
         );
  OAI22XL U1947 ( .A0(n618), .A1(n575), .B0(n334), .B1(n233), .Y(\C2/Z_9 ) );
  AOI222XL U1948 ( .A0(n574), .A1(n355), .B0(n616), .B1(n109), .C0(n632), .C1(
        read_cntr[1]), .Y(n575) );
  OAI22XL U1949 ( .A0(n618), .A1(n573), .B0(n334), .B1(n284), .Y(\C2/Z_10 ) );
  AO22X1 U1950 ( .A0(n610), .A1(n112), .B0(n616), .B1(n110), .Y(n570) );
  AO21X1 U1951 ( .A0(curr_photo_addr[11]), .A1(n338), .B0(si_sel), .Y(
        \C1/Z_11 ) );
  OAI22XL U1952 ( .A0(n618), .A1(n569), .B0(n334), .B1(n250), .Y(\C2/Z_11 ) );
  AO22X1 U1953 ( .A0(n610), .A1(n109), .B0(n616), .B1(write_addr[11]), .Y(n567) );
  OAI22XL U1954 ( .A0(n618), .A1(n566), .B0(n334), .B1(n244), .Y(\C2/Z_12 ) );
  OAI2BB2XL U1955 ( .B0(n275), .B1(n594), .A0N(n610), .A1N(n110), .Y(n564) );
  AO21X1 U1956 ( .A0(n2131), .A1(n659), .B0(n2130), .Y(n572) );
  AO21X1 U1957 ( .A0(curr_photo_addr[13]), .A1(n338), .B0(si_sel), .Y(
        \C1/Z_13 ) );
  OAI22XL U1958 ( .A0(n618), .A1(n562), .B0(n334), .B1(n317), .Y(\C2/Z_13 ) );
  AO22X1 U1959 ( .A0(n610), .A1(write_addr[11]), .B0(n616), .B1(write_addr[13]), .Y(n559) );
  AO21X1 U1960 ( .A0(curr_photo_addr[14]), .A1(n338), .B0(si_sel), .Y(
        \C1/Z_14 ) );
  OAI22XL U1961 ( .A0(n618), .A1(n557), .B0(n334), .B1(n243), .Y(\C2/Z_14 ) );
  OAI22XL U1962 ( .A0(n608), .A1(n554), .B0(n594), .B1(n274), .Y(n555) );
  AO21X1 U1963 ( .A0(curr_photo_addr[15]), .A1(n338), .B0(si_sel), .Y(
        \C1/Z_15 ) );
  OAI22XL U1964 ( .A0(n618), .A1(n553), .B0(n334), .B1(n319), .Y(\C2/Z_15 ) );
  OAI22XL U1965 ( .A0(n608), .A1(n550), .B0(n594), .B1(n2203), .Y(n551) );
  OAI22XL U1966 ( .A0(n618), .A1(n549), .B0(n334), .B1(n225), .Y(\C2/Z_16 ) );
  OAI22XL U1967 ( .A0(n2231), .A1(n608), .B0(n594), .B1(n2230), .Y(n547) );
  OA21XL U1968 ( .A0(n2201), .A1(write_addr[14]), .B0(n2202), .Y(n419) );
  OAI22XL U1969 ( .A0(n618), .A1(n546), .B0(n334), .B1(n320), .Y(\C2/Z_17 ) );
  OAI22XL U1970 ( .A0(n2232), .A1(n608), .B0(n594), .B1(n318), .Y(n544) );
  OAI22XL U1971 ( .A0(n618), .A1(n543), .B0(n334), .B1(n247), .Y(\C2/Z_18 ) );
  AO22X1 U1972 ( .A0(n355), .A1(n540), .B0(n616), .B1(write_addr[18]), .Y(n541) );
  OA21XL U1973 ( .A0(global_cntr[15]), .A1(n370), .B0(n668), .Y(n642) );
  OA21XL U1974 ( .A0(global_cntr[13]), .A1(n368), .B0(n369), .Y(n644) );
  OA21XL U1975 ( .A0(global_cntr[4]), .A1(n361), .B0(n362), .Y(n654) );
  AOI2BB1X1 U1976 ( .A0N(global_cntr[3]), .A1N(n656), .B0(n361), .Y(n655) );
  NOR2X1 U1977 ( .A(n375), .B(n374), .Y(n638) );
  NOR2X1 U1978 ( .A(n375), .B(n371), .Y(n640) );
  NAND2XL U1979 ( .A(n257), .B(n1189), .Y(n1190) );
  OAI2BB1X1 U1980 ( .A0N(n1070), .A1N(n1071), .B0(n398), .Y(n622) );
  OR2X1 U1981 ( .A(n735), .B(n1449), .Y(n219) );
  OA21XL U1982 ( .A0(n733), .A1(n219), .B0(n732), .Y(n242) );
  OR2X1 U1983 ( .A(global_cntr[8]), .B(global_cntr[11]), .Y(n926) );
  AO21X1 U1984 ( .A0(n233), .A1(n673), .B0(n648), .Y(n667) );
  OAI21XL U1985 ( .A0(n651), .A1(next_glb_cntr[6]), .B0(n650), .Y(n666) );
  OR4X1 U1986 ( .A(n645), .B(n644), .C(n643), .D(n642), .Y(n674) );
  OAI31XL U1987 ( .A0(n111), .A1(write_cntr[5]), .A2(write_cntr[6]), .B0(
        write_cntr[9]), .Y(n680) );
  OAI21XL U1988 ( .A0(n245), .A1(n680), .B0(n221), .Y(n681) );
  OA22X1 U1989 ( .A0(n2218), .A1(n687), .B0(n661), .B1(n1435), .Y(n685) );
  OAI21XL U1990 ( .A0(n714), .A1(n723), .B0(n245), .Y(n715) );
  NAND3BX1 U1991 ( .AN(n908), .B(n1977), .C(n180), .Y(n902) );
  OAI21XL U1992 ( .A0(n219), .A1(n735), .B0(n1449), .Y(n734) );
  OAI21XL U1993 ( .A0(n742), .A1(n737), .B0(n740), .Y(n738) );
  OAI21XL U1994 ( .A0(n744), .A1(n2135), .B0(n743), .Y(n741) );
  OAI21XL U1995 ( .A0(n2135), .A1(n746), .B0(n747), .Y(n745) );
  OAI21XL U1996 ( .A0(n759), .A1(n756), .B0(n758), .Y(n757) );
  OAI21XL U1997 ( .A0(n764), .A1(n2145), .B0(n763), .Y(n762) );
  OAI21XL U1998 ( .A0(n180), .A1(n765), .B0(n768), .Y(n766) );
  OAI21XL U1999 ( .A0(n2145), .A1(n770), .B0(n771), .Y(n769) );
  NAND3BX1 U2000 ( .AN(n776), .B(n775), .C(n1978), .Y(n773) );
  OAI21XL U2001 ( .A0(n779), .A1(n776), .B0(n778), .Y(n777) );
  AOI2BB2X1 U2002 ( .B0(n1997), .B1(n2157), .A0N(n1997), .A1N(n2157), .Y(n796)
         );
  AOI2BB2X1 U2003 ( .B0(n2164), .B1(n2017), .A0N(n2164), .A1N(n2017), .Y(n809)
         );
  OAI2BB1X1 U2004 ( .A0N(n801), .A1N(n800), .B0(n799), .Y(n802) );
  AOI2BB2X1 U2005 ( .B0(n2021), .B1(n2170), .A0N(n2021), .A1N(n2170), .Y(n824)
         );
  OAI2BB1X1 U2006 ( .A0N(n819), .A1N(n823), .B0(n164), .Y(n820) );
  OAI21XL U2007 ( .A0(n2119), .A1(n833), .B0(n834), .Y(n832) );
  AO21X1 U2008 ( .A0(n840), .A1(n839), .B0(n838), .Y(n841) );
  AOI2BB2X1 U2009 ( .B0(n1442), .B1(n2124), .A0N(n1442), .A1N(n2124), .Y(n2052) );
  OR2X1 U2010 ( .A(n1442), .B(n850), .Y(n848) );
  OAI22XL U2011 ( .A0(n2042), .A1(n853), .B0(n852), .B1(n2041), .Y(n854) );
  AOI2BB1X1 U2012 ( .A0N(work_cntr[4]), .A1N(n898), .B0(n887), .Y(n1747) );
  AO21X1 U2013 ( .A0(n261), .A1(n885), .B0(n888), .Y(n1718) );
  OAI2BB1X1 U2014 ( .A0N(n263), .A1N(n886), .B0(n885), .Y(n1731) );
  AO21X1 U2015 ( .A0(n268), .A1(n893), .B0(n894), .Y(n1658) );
  NAND3BX1 U2016 ( .AN(n895), .B(work_cntr[16]), .C(work_cntr[15]), .Y(n1627)
         );
  AO21X1 U2017 ( .A0(n222), .A1(n1627), .B0(n148), .Y(n1618) );
  OAI21XL U2018 ( .A0(n1955), .A1(n286), .B0(n914), .Y(n913) );
  OR4X1 U2019 ( .A(n107), .B(global_cntr[5]), .C(global_cntr[9]), .D(
        global_cntr[14]), .Y(n925) );
  OAI22XL U2020 ( .A0(work_cntr[17]), .A1(n1792), .B0(n222), .B1(n259), .Y(
        n934) );
  AOI2BB2X1 U2021 ( .B0(n260), .B1(n939), .A0N(n260), .A1N(n939), .Y(n946) );
  OAI21XL U2022 ( .A0(n958), .A1(work_cntr[13]), .B0(n957), .Y(n956) );
  AO21X1 U2023 ( .A0(n980), .A1(n975), .B0(work_cntr[11]), .Y(n977) );
  OAI21XL U2024 ( .A0(n975), .A1(work_cntr[11]), .B0(n974), .Y(n973) );
  OAI21XL U2025 ( .A0(n986), .A1(work_cntr[10]), .B0(n989), .Y(n987) );
  AO21X1 U2026 ( .A0(n1008), .A1(n1001), .B0(work_cntr[8]), .Y(n1003) );
  OAI21XL U2027 ( .A0(n1001), .A1(work_cntr[8]), .B0(n1004), .Y(n1002) );
  OR2X1 U2028 ( .A(n1012), .B(n1006), .Y(n1013) );
  AO21X1 U2029 ( .A0(n1013), .A1(n1011), .B0(work_cntr[7]), .Y(n1014) );
  OAI21XL U2030 ( .A0(n1011), .A1(work_cntr[7]), .B0(n1010), .Y(n1009) );
  OR2X1 U2031 ( .A(n1017), .B(n1016), .Y(n1024) );
  AO21X1 U2032 ( .A0(n1024), .A1(n1021), .B0(work_cntr[6]), .Y(n1018) );
  OA21XL U2033 ( .A0(n263), .A1(n1023), .B0(n1018), .Y(n1026) );
  AO21X1 U2034 ( .A0(n1029), .A1(n1027), .B0(work_cntr[5]), .Y(n1030) );
  OAI21XL U2035 ( .A0(n1027), .A1(work_cntr[5]), .B0(n1026), .Y(n1025) );
  OR2X1 U2036 ( .A(n1033), .B(n160), .Y(n1041) );
  AO21X1 U2037 ( .A0(n1041), .A1(n1035), .B0(work_cntr[4]), .Y(n1037) );
  OAI21XL U2038 ( .A0(n1035), .A1(work_cntr[4]), .B0(n1038), .Y(n1036) );
  OAI21XL U2039 ( .A0(n1046), .A1(N1184), .B0(n1048), .Y(n1047) );
  OAI21XL U2040 ( .A0(n1057), .A1(N1183), .B0(n1060), .Y(n1058) );
  OR2X1 U2041 ( .A(n1320), .B(work_cntr[13]), .Y(n1301) );
  AO21X1 U2042 ( .A0(n1090), .A1(n215), .B0(n1074), .Y(n1112) );
  OR2X1 U2043 ( .A(n1080), .B(n1082), .Y(n1083) );
  AOI222XL U2044 ( .A0(n1092), .A1(n1089), .B0(n1092), .B1(work_cntr[16]), 
        .C0(n1089), .C1(n211), .Y(n1087) );
  AOI2BB2X1 U2045 ( .B0(n1088), .B1(n1087), .A0N(n1088), .A1N(n1086), .Y(n1098) );
  OR2X1 U2046 ( .A(n1092), .B(n211), .Y(n1097) );
  OAI21XL U2047 ( .A0(n1095), .A1(n1094), .B0(n211), .Y(n1096) );
  OAI21XL U2048 ( .A0(work_cntr[15]), .A1(n1112), .B0(n1098), .Y(n1100) );
  OAI21XL U2049 ( .A0(n215), .A1(n1114), .B0(n1111), .Y(n1102) );
  NOR3BXL U2050 ( .AN(n1112), .B(n1111), .C(n1109), .Y(n1105) );
  NAND3BX1 U2051 ( .AN(n1105), .B(n1106), .C(n1114), .Y(n1122) );
  OAI21XL U2052 ( .A0(n1109), .A1(n1111), .B0(n1112), .Y(n1110) );
  OAI21XL U2053 ( .A0(work_cntr[13]), .A1(n1126), .B0(n1113), .Y(n1116) );
  AOI2BB2X1 U2054 ( .B0(n1117), .B1(n1116), .A0N(n1117), .A1N(n1115), .Y(n1121) );
  OAI21XL U2055 ( .A0(work_cntr[12]), .A1(n1129), .B0(n1121), .Y(n1118) );
  AOI2BB2X1 U2056 ( .B0(work_cntr[10]), .B1(n1124), .A0N(work_cntr[10]), .A1N(
        n1124), .Y(n1135) );
  OAI21XL U2057 ( .A0(work_cntr[11]), .A1(n1142), .B0(n1128), .Y(n1131) );
  AO22X1 U2058 ( .A0(n1132), .A1(n1131), .B0(n1130), .B1(n1129), .Y(n1143) );
  OAI21XL U2059 ( .A0(work_cntr[10]), .A1(n204), .B0(n1133), .Y(n1134) );
  AOI2BB2X1 U2060 ( .B0(n1136), .B1(n1135), .A0N(n1136), .A1N(n1134), .Y(n1144) );
  AOI2BB1X1 U2061 ( .A0N(n1139), .A1N(n262), .B0(n1138), .Y(n1149) );
  AOI2BB2X1 U2062 ( .B0(work_cntr[7]), .B1(n1140), .A0N(work_cntr[7]), .A1N(
        n1140), .Y(n1151) );
  AO21X1 U2063 ( .A0(n262), .A1(n1160), .B0(n1156), .Y(n1147) );
  AOI2BB2X1 U2064 ( .B0(n1148), .B1(n1149), .A0N(n1148), .A1N(n1147), .Y(n1157) );
  OA21XL U2065 ( .A0(n1156), .A1(n1155), .B0(n1154), .Y(n1161) );
  OAI21XL U2066 ( .A0(work_cntr[7]), .A1(n1169), .B0(n1158), .Y(n1159) );
  AO21X1 U2067 ( .A0(n263), .A1(n1175), .B0(n1170), .Y(n1162) );
  OA21XL U2068 ( .A0(n1170), .A1(n1169), .B0(n1168), .Y(n1176) );
  OAI21XL U2069 ( .A0(work_cntr[5]), .A1(n1182), .B0(n1173), .Y(n1174) );
  AO21X1 U2070 ( .A0(n1180), .A1(n1183), .B0(n1177), .Y(n1178) );
  AOI221XL U2071 ( .A0(n1766), .A1(n1185), .B0(n1184), .B1(n1758), .C0(n1187), 
        .Y(n1186) );
  AO21X1 U2072 ( .A0(n257), .A1(n1783), .B0(n1197), .Y(n1194) );
  AOI2BB2X1 U2073 ( .B0(n1188), .B1(n1756), .A0N(n1188), .A1N(n1187), .Y(n1192) );
  AOI2BB2X1 U2074 ( .B0(n1778), .B1(n1195), .A0N(n1778), .A1N(n1195), .Y(n2223) );
  OR2X1 U2075 ( .A(n1203), .B(n1278), .Y(n1206) );
  AOI2BB2X1 U2076 ( .B0(n248), .B1(n1205), .A0N(n248), .A1N(n1205), .Y(n1211)
         );
  AOI2BB2X1 U2077 ( .B0(write_cntr[12]), .B1(n1206), .A0N(write_cntr[12]), 
        .A1N(n1206), .Y(n1209) );
  NAND3BX1 U2078 ( .AN(n221), .B(write_cntr[8]), .C(n1223), .Y(n1207) );
  NAND3BX1 U2079 ( .AN(n166), .B(n1209), .C(n1207), .Y(n1216) );
  AOI2BB2X1 U2080 ( .B0(n166), .B1(n1210), .A0N(n166), .A1N(n1210), .Y(n1226)
         );
  AOI2BB2X1 U2081 ( .B0(n1219), .B1(n1218), .A0N(n1219), .A1N(n1217), .Y(n1230) );
  NAND3BX1 U2082 ( .AN(n1241), .B(n1233), .C(n1243), .Y(n1244) );
  AOI2BB2X1 U2083 ( .B0(n1232), .B1(n1231), .A0N(n1232), .A1N(n1230), .Y(n1245) );
  AOI2BB2X1 U2084 ( .B0(n1241), .B1(n1240), .A0N(n1241), .A1N(n1240), .Y(n1253) );
  OAI21XL U2085 ( .A0(n1251), .A1(n1248), .B0(n1250), .Y(n1247) );
  AOI2BB2X1 U2086 ( .B0(n1259), .B1(n1258), .A0N(n1259), .A1N(n1258), .Y(n1262) );
  AOI2BB2X1 U2087 ( .B0(n1261), .B1(n1260), .A0N(n1261), .A1N(n1260), .Y(n1271) );
  OAI21XL U2088 ( .A0(write_cntr[4]), .A1(n1440), .B0(write_cntr[3]), .Y(n1265) );
  OAI221XL U2089 ( .A0(n1268), .A1(n1265), .B0(n1269), .B1(n1268), .C0(n1267), 
        .Y(n1266) );
  OAI31XL U2090 ( .A0(n1269), .A1(n1268), .A2(n1267), .B0(n1266), .Y(n1270) );
  OA21XL U2091 ( .A0(n1274), .A1(n1275), .B0(n1270), .Y(n1273) );
  OAI21XL U2092 ( .A0(n227), .A1(N76), .B0(n1414), .Y(n1284) );
  OAI2BB1X1 U2093 ( .A0N(n1790), .A1N(work_cntr[16]), .B0(n1289), .Y(n1292) );
  OA21XL U2094 ( .A0(n1293), .A1(n1292), .B0(n1298), .Y(n1296) );
  AOI2BB2X1 U2095 ( .B0(n1304), .B1(n1303), .A0N(n1304), .A1N(n1302), .Y(n1307) );
  AOI2BB1X1 U2096 ( .A0N(n1307), .A1N(n1311), .B0(n1306), .Y(n1309) );
  OR2X1 U2097 ( .A(n1323), .B(n1325), .Y(n1313) );
  OR2X1 U2098 ( .A(n1314), .B(n1313), .Y(n1310) );
  OAI2BB1X1 U2099 ( .A0N(n1335), .A1N(n1333), .B0(n1324), .Y(n1330) );
  AOI2BB2X1 U2100 ( .B0(n1331), .B1(n1330), .A0N(n1331), .A1N(n1329), .Y(n1336) );
  AOI2BB2X1 U2101 ( .B0(n1335), .B1(n1334), .A0N(n1335), .A1N(n1334), .Y(n1339) );
  AOI2BB2X1 U2102 ( .B0(work_cntr[11]), .B1(n1808), .A0N(work_cntr[11]), .A1N(
        n1808), .Y(n1340) );
  AOI2BB2X1 U2103 ( .B0(n1342), .B1(n1341), .A0N(n1342), .A1N(n1341), .Y(n1343) );
  OAI21XL U2104 ( .A0(n1350), .A1(n1346), .B0(n1343), .Y(n1344) );
  OAI21XL U2105 ( .A0(n1351), .A1(n1349), .B0(n1350), .Y(n1348) );
  NAND3BX1 U2106 ( .AN(n175), .B(n1369), .C(n1363), .Y(n1370) );
  AOI2BB2X1 U2107 ( .B0(n1366), .B1(n1359), .A0N(n1366), .A1N(n1359), .Y(n1361) );
  OAI21XL U2108 ( .A0(n1369), .A1(n1368), .B0(n1367), .Y(n1371) );
  AOI2BB2X1 U2109 ( .B0(n1375), .B1(n1374), .A0N(n1375), .A1N(n1374), .Y(n1395) );
  AOI2BB2X1 U2110 ( .B0(n1379), .B1(n175), .A0N(n1379), .A1N(n175), .Y(n1381)
         );
  NAND3BX1 U2111 ( .AN(n1384), .B(n1395), .C(n1386), .Y(n1388) );
  AOI2BB2X1 U2112 ( .B0(n1387), .B1(n1386), .A0N(n1387), .A1N(n1386), .Y(n1389) );
  AOI221XL U2113 ( .A0(work_cntr[4]), .A1(n229), .B0(n1396), .B1(work_cntr[5]), 
        .C0(n1401), .Y(n1393) );
  AOI2BB2X1 U2114 ( .B0(n223), .B1(n1398), .A0N(n223), .A1N(n1398), .Y(n1408)
         );
  OAI21XL U2115 ( .A0(n1402), .A1(n1400), .B0(n1401), .Y(n1399) );
  AOI2BB2X1 U2116 ( .B0(n1405), .B1(n1404), .A0N(n1405), .A1N(n1404), .Y(n1407) );
  AOI2BB1X1 U2117 ( .A0N(n1411), .A1N(n1407), .B0(n1406), .Y(n1421) );
  OAI22XL U2118 ( .A0(N1182), .A1(N1183), .B0(n1911), .B1(n1421), .Y(n1409) );
  OAI21XL U2119 ( .A0(n1783), .A1(n1414), .B0(n1413), .Y(n1415) );
  AOI2BB2X1 U2120 ( .B0(n1432), .B1(n1429), .A0N(n1417), .A1N(n1426), .Y(n1418) );
  ADDFXL U2121 ( .A(N1183), .B(n1421), .CI(n1420), .CO(n1424), .S(n1432) );
  OAI21XL U2122 ( .A0(n1425), .A1(n1423), .B0(n1424), .Y(n1422) );
  NOR2X1 U2123 ( .A(n1430), .B(n2241), .Y(expand_sel[3]) );
  OAI2BB2XL U2124 ( .B0(n1443), .B1(im_wen_n), .A0N(write_cntr[2]), .A1N(n147), 
        .Y(n353) );
  AO22X1 U2125 ( .A0(n147), .A1(write_cntr[0]), .B0(n360), .B1(n2050), .Y(n349) );
  OAI2BB2XL U2126 ( .B0(n2004), .B1(im_wen_n), .A0N(write_cntr[6]), .A1N(n147), 
        .Y(n346) );
  AOI2BB2X1 U2127 ( .B0(n235), .B1(im_wen_n), .A0N(n1448), .A1N(n147), .Y(n341) );
  AOI2BB2X1 U2128 ( .B0(next_work_cntr[17]), .B1(n1461), .A0N(
        next_work_cntr[17]), .A1N(n1461), .Y(n1476) );
  OA21XL U2129 ( .A0(n173), .A1(n1472), .B0(n1468), .Y(n1465) );
  AOI2BB2X1 U2130 ( .B0(n1478), .B1(n1477), .A0N(n1478), .A1N(n1476), .Y(n1481) );
  OAI2BB2XL U2131 ( .B0(n1489), .B1(n1488), .A0N(n1489), .A1N(n1488), .Y(n1491) );
  AOI2BB2X1 U2132 ( .B0(n1499), .B1(next_work_cntr[11]), .A0N(n1499), .A1N(
        next_work_cntr[11]), .Y(n1517) );
  OAI21XL U2133 ( .A0(n1515), .A1(n1513), .B0(n1514), .Y(n1512) );
  AOI2BB2X1 U2134 ( .B0(n1522), .B1(n1518), .A0N(n1522), .A1N(n1518), .Y(n1527) );
  AO21X1 U2135 ( .A0(n1537), .A1(n1547), .B0(n1548), .Y(n1549) );
  AOI2BB2X1 U2136 ( .B0(n1541), .B1(n1540), .A0N(n1541), .A1N(n1540), .Y(n1554) );
  OAI21XL U2137 ( .A0(n1549), .A1(n1546), .B0(n1556), .Y(n1559) );
  OAI21XL U2138 ( .A0(n1563), .A1(n1562), .B0(n1551), .Y(n1552) );
  NAND3BX1 U2139 ( .AN(n1575), .B(n1574), .C(n1571), .Y(n1564) );
  OAI21XL U2140 ( .A0(n1574), .A1(n1571), .B0(n1564), .Y(n1565) );
  OA21XL U2141 ( .A0(n1568), .A1(n1567), .B0(n1566), .Y(n1582) );
  AOI2BB2X1 U2142 ( .B0(n1583), .B1(n1584), .A0N(n1583), .A1N(n1584), .Y(n1601) );
  OAI21XL U2143 ( .A0(n1591), .A1(n1589), .B0(n1590), .Y(n1588) );
  AOI2BB2X1 U2144 ( .B0(n1594), .B1(n1593), .A0N(n1594), .A1N(n1593), .Y(n1607) );
  OAI22XL U2145 ( .A0(n1597), .A1(n1598), .B0(next_work_cntr[19]), .B1(n1596), 
        .Y(n1605) );
  OAI21XL U2146 ( .A0(n1603), .A1(n1601), .B0(n1600), .Y(n1602) );
  OAI21XL U2147 ( .A0(n1603), .A1(n1606), .B0(n1602), .Y(n1604) );
  OAI21XL U2148 ( .A0(n1610), .A1(n1609), .B0(n1608), .Y(n1611) );
  OAI21XL U2149 ( .A0(n1613), .A1(n1612), .B0(n1611), .Y(n1617) );
  OAI21XL U2150 ( .A0(n656), .A1(n1615), .B0(n1614), .Y(n1616) );
  OA22X1 U2151 ( .A0(n259), .A1(n1623), .B0(n1622), .B1(n1621), .Y(n1630) );
  AO22X1 U2152 ( .A0(n1627), .A1(n1626), .B0(n1798), .B1(n148), .Y(n1631) );
  NAND3BX1 U2153 ( .AN(n1629), .B(n1631), .C(n1633), .Y(n1628) );
  OAI2BB1X1 U2154 ( .A0N(n1629), .A1N(n1632), .B0(n1628), .Y(n1636) );
  AO21X1 U2155 ( .A0(n1637), .A1(n1641), .B0(n1640), .Y(n1643) );
  OAI21XL U2156 ( .A0(n1641), .A1(n1640), .B0(n1644), .Y(n1642) );
  OR2X1 U2157 ( .A(n1650), .B(n1645), .Y(n1654) );
  AO21X1 U2158 ( .A0(n1654), .A1(n1649), .B0(n1648), .Y(n1651) );
  OA21XL U2159 ( .A0(n1652), .A1(n1653), .B0(n1651), .Y(n1663) );
  AO21X1 U2160 ( .A0(n1656), .A1(n1660), .B0(n1659), .Y(n1662) );
  OAI21XL U2161 ( .A0(n1660), .A1(n1659), .B0(n1663), .Y(n1661) );
  OR2X1 U2162 ( .A(n156), .B(n1664), .Y(n1674) );
  AO21X1 U2163 ( .A0(n1674), .A1(n1668), .B0(n1667), .Y(n1670) );
  OA21XL U2164 ( .A0(n1671), .A1(n1673), .B0(n1670), .Y(n1683) );
  AO21X1 U2165 ( .A0(n1676), .A1(n1680), .B0(n1679), .Y(n1682) );
  OAI21XL U2166 ( .A0(n1680), .A1(n1679), .B0(n1683), .Y(n1681) );
  OR2X1 U2167 ( .A(n157), .B(n1684), .Y(n1694) );
  AO21X1 U2168 ( .A0(n1694), .A1(n1688), .B0(n1687), .Y(n1690) );
  OA21XL U2169 ( .A0(n1691), .A1(n1693), .B0(n1690), .Y(n1703) );
  AO21X1 U2170 ( .A0(n1696), .A1(n1700), .B0(n1699), .Y(n1702) );
  OAI21XL U2171 ( .A0(n1700), .A1(n1699), .B0(n1703), .Y(n1701) );
  OR2X1 U2172 ( .A(n158), .B(n1704), .Y(n1714) );
  AO21X1 U2173 ( .A0(n1714), .A1(n1708), .B0(n1707), .Y(n1710) );
  OA21XL U2174 ( .A0(n1711), .A1(n1713), .B0(n1710), .Y(n1723) );
  AO21X1 U2175 ( .A0(n1716), .A1(n1720), .B0(n1719), .Y(n1722) );
  OAI21XL U2176 ( .A0(n1720), .A1(n1719), .B0(n1723), .Y(n1721) );
  OR2X1 U2177 ( .A(n159), .B(n1724), .Y(n1734) );
  AO21X1 U2178 ( .A0(n1734), .A1(n1728), .B0(n1727), .Y(n1730) );
  AO21X1 U2179 ( .A0(n1736), .A1(n1740), .B0(n1739), .Y(n1742) );
  OAI21XL U2180 ( .A0(n1740), .A1(n1739), .B0(n152), .Y(n1741) );
  OR2X1 U2181 ( .A(n1744), .B(n1749), .Y(n1750) );
  AO21X1 U2182 ( .A0(n1750), .A1(n1748), .B0(n1747), .Y(n1751) );
  OAI31XL U2183 ( .A0(n1748), .A1(n1747), .A2(n1746), .B0(n1745), .Y(n1755) );
  OA21XL U2184 ( .A0(n1753), .A1(n1752), .B0(n1751), .Y(n1762) );
  AO21X1 U2185 ( .A0(n1765), .A1(n1759), .B0(n1758), .Y(n1761) );
  OAI21XL U2186 ( .A0(n1759), .A1(n1758), .B0(n1762), .Y(n1760) );
  OR2X1 U2187 ( .A(n1763), .B(n161), .Y(n1771) );
  AO21X1 U2188 ( .A0(n1771), .A1(n1769), .B0(n1766), .Y(n1772) );
  OAI21XL U2189 ( .A0(n1769), .A1(n1766), .B0(n1768), .Y(n1767) );
  OA21XL U2190 ( .A0(n1779), .A1(n1778), .B0(n1780), .Y(n1787) );
  OAI31XL U2191 ( .A0(n1784), .A1(n1783), .A2(n1782), .B0(n1781), .Y(n1785) );
  AOI2BB1X1 U2192 ( .A0N(n1789), .A1N(n258), .B0(n1785), .Y(n1786) );
  AOI2BB2X1 U2193 ( .B0(n222), .B1(n1802), .A0N(n222), .A1N(n1802), .Y(n1799)
         );
  OA21XL U2194 ( .A0(n1793), .A1(n1792), .B0(n1799), .Y(n1797) );
  AOI2BB2X1 U2195 ( .B0(n1795), .B1(n1894), .A0N(n1794), .A1N(n236), .Y(n1796)
         );
  OAI2BB2XL U2196 ( .B0(n1804), .B1(n260), .A0N(n1822), .A1N(n1814), .Y(n1806)
         );
  AOI2BB2X1 U2197 ( .B0(n214), .B1(n1816), .A0N(n214), .A1N(n1816), .Y(n1820)
         );
  AO21X1 U2198 ( .A0(n264), .A1(n1825), .B0(n214), .Y(n1817) );
  AOI2BB2X1 U2199 ( .B0(n1818), .B1(n1817), .A0N(n1818), .A1N(n1816), .Y(n1829) );
  OAI21XL U2200 ( .A0(n215), .A1(n1835), .B0(n1829), .Y(n1819) );
  AOI2BB2X1 U2201 ( .B0(n1820), .B1(n1825), .A0N(n1820), .A1N(n1819), .Y(n1831) );
  AO21X1 U2202 ( .A0(n1827), .A1(n1826), .B0(n1825), .Y(n1828) );
  OAI21XL U2203 ( .A0(work_cntr[13]), .A1(n1850), .B0(n1832), .Y(n1833) );
  AO22X1 U2204 ( .A0(n1836), .A1(n1835), .B0(n1834), .B1(n1833), .Y(n1851) );
  AO21X1 U2205 ( .A0(n209), .A1(n1854), .B0(n1851), .Y(n1837) );
  AO21X1 U2206 ( .A0(work_cntr[10]), .A1(n1845), .B0(n1844), .Y(n1867) );
  OAI21XL U2207 ( .A0(work_cntr[11]), .A1(n1867), .B0(n1852), .Y(n1853) );
  AOI2BB2X1 U2208 ( .B0(n1855), .B1(n1854), .A0N(n1855), .A1N(n1853), .Y(n1868) );
  OAI21XL U2209 ( .A0(work_cntr[10]), .A1(n1870), .B0(n1860), .Y(n1857) );
  OAI21XL U2210 ( .A0(work_cntr[9]), .A1(n1880), .B0(n1869), .Y(n1872) );
  AO22X1 U2211 ( .A0(n1873), .A1(n1872), .B0(n1871), .B1(n1870), .Y(n1881) );
  OAI21XL U2212 ( .A0(work_cntr[8]), .A1(n1888), .B0(n1874), .Y(n1875) );
  AOI2BB2X1 U2213 ( .B0(n1877), .B1(n1876), .A0N(n1877), .A1N(n1875), .Y(n1889) );
  AO21X1 U2214 ( .A0(n261), .A1(n1898), .B0(n1889), .Y(n1882) );
  AOI2BB2X1 U2215 ( .B0(n1884), .B1(n1883), .A0N(n1884), .A1N(n1882), .Y(n1897) );
  OAI21XL U2216 ( .A0(work_cntr[6]), .A1(n178), .B0(n1890), .Y(n1891) );
  AO21X1 U2217 ( .A0(n229), .A1(n1915), .B0(n1903), .Y(n1899) );
  NAND3BX1 U2218 ( .AN(n1904), .B(n1903), .C(n178), .Y(n1905) );
  OAI21XL U2219 ( .A0(work_cntr[4]), .A1(n1919), .B0(n1908), .Y(n1906) );
  AOI2BB2X1 U2220 ( .B0(n1907), .B1(n1915), .A0N(n1907), .A1N(n1906), .Y(n1910) );
  AOI2BB2X1 U2221 ( .B0(N1183), .B1(n1925), .A0N(N1183), .A1N(n1925), .Y(n1927) );
  OAI2BB1X1 U2222 ( .A0N(n1929), .A1N(N1182), .B0(n258), .Y(n1926) );
  OAI21XL U2223 ( .A0(n1929), .A1(N1182), .B0(n1928), .Y(n1930) );
  AOI2BB2X1 U2224 ( .B0(n1931), .B1(n2237), .A0N(n1931), .A1N(n1930), .Y(n1932) );
  AO22X1 U2225 ( .A0(cr_read_cntr[4]), .A1(n1945), .B0(n322), .B1(n1949), .Y(
        n312) );
  OAI22XL U2226 ( .A0(cr_read_cntr[6]), .A1(n1950), .B0(n286), .B1(n1952), .Y(
        n310) );
  OA21XL U2227 ( .A0(cr_read_cntr[7]), .A1(n1954), .B0(n1953), .Y(n309) );
  AO22X1 U2228 ( .A0(n1955), .A1(n1954), .B0(cr_read_cntr[8]), .B1(n1953), .Y(
        n308) );
  AOI2BB2X1 U2229 ( .B0(n1956), .B1(write_addr[17]), .A0N(n1956), .A1N(
        write_addr[17]), .Y(n2210) );
  AOI2BB2X1 U2230 ( .B0(n1957), .B1(write_addr[16]), .A0N(n1957), .A1N(
        write_addr[16]), .Y(n2207) );
  AO21X1 U2231 ( .A0(n1959), .A1(n275), .B0(n1960), .Y(n2188) );
  AOI2BB2X1 U2232 ( .B0(n2066), .B1(n238), .A0N(n2066), .A1N(n238), .Y(n2075)
         );
  OAI21XL U2233 ( .A0(n112), .A1(n2045), .B0(n1974), .Y(n1970) );
  AO21X1 U2234 ( .A0(n2083), .A1(n2002), .B0(n2018), .Y(n2019) );
  AOI2BB2X1 U2235 ( .B0(n2004), .B1(n2088), .A0N(n2003), .A1N(n2018), .Y(n2005) );
  AOI2BB2X1 U2236 ( .B0(n2006), .B1(n2005), .A0N(n2006), .A1N(n2005), .Y(n2030) );
  AOI2BB2X1 U2237 ( .B0(n2009), .B1(n2007), .A0N(n2009), .A1N(n2007), .Y(n2032) );
  OA21XL U2238 ( .A0(n2016), .A1(n2015), .B0(n2014), .Y(n2036) );
  OAI22XL U2239 ( .A0(n2030), .A1(n2031), .B0(n2028), .B1(n2027), .Y(n2029) );
  OAI2BB1X1 U2240 ( .A0N(n2031), .A1N(n2030), .B0(n2029), .Y(n2033) );
  OAI21XL U2241 ( .A0(n2036), .A1(n2035), .B0(n2034), .Y(n2037) );
  AOI2BB2X1 U2242 ( .B0(n2040), .B1(n2039), .A0N(n2040), .A1N(n2039), .Y(n2071) );
  OAI21XL U2243 ( .A0(n2046), .A1(n2045), .B0(n2044), .Y(n2047) );
  OR2X1 U2244 ( .A(n2059), .B(n2050), .Y(n2051) );
  OR2X1 U2245 ( .A(n2059), .B(n2058), .Y(n2070) );
  OAI221XL U2246 ( .A0(n2062), .A1(n2061), .B0(n2060), .B1(n2061), .C0(n2070), 
        .Y(n2063) );
  AOI2BB2X1 U2247 ( .B0(n2074), .B1(n2073), .A0N(n2074), .A1N(n2073), .Y(n2065) );
  AOI2BB2X1 U2248 ( .B0(n2077), .B1(n2065), .A0N(n2077), .A1N(n2065), .Y(n2067) );
  AO21X1 U2249 ( .A0(n2071), .A1(n2070), .B0(n2069), .Y(n2072) );
  AOI222XL U2250 ( .A0(n2077), .A1(n2074), .B0(n2077), .B1(n2073), .C0(n2074), 
        .C1(n2073), .Y(\intadd_3/CI ) );
  ADDFXL U2251 ( .A(n2078), .B(n2077), .CI(n2076), .CO(n2079), .S(n2068) );
  ADDFXL U2252 ( .A(n2086), .B(n2085), .CI(n2084), .CO(\intadd_3/B[2] ), .S(
        \intadd_3/A[1] ) );
  OAI21XL U2253 ( .A0(n2098), .A1(\intadd_3/n1 ), .B0(n659), .Y(n2089) );
  ADDFXL U2254 ( .A(n2095), .B(n2094), .CI(n2093), .CO(n2096), .S(
        \intadd_3/A[2] ) );
  OAI21XL U2255 ( .A0(n2110), .A1(n2109), .B0(n2108), .Y(n2114) );
  ADDFXL U2256 ( .A(next_cr_x[5]), .B(n2111), .CI(n2107), .CO(n2112), .S(n2100) );
  AOI2BB2X1 U2257 ( .B0(\DP_OP_436J1_125_1438/n25 ), .B1(n2122), .A0N(
        \DP_OP_436J1_125_1438/n25 ), .A1N(n2122), .Y(n2117) );
  ADDFXL U2258 ( .A(n251), .B(next_cr_x[6]), .CI(n2124), .CO(n2132), .S(n2121)
         );
  AOI2BB2X1 U2259 ( .B0(n237), .B1(n2138), .A0N(n237), .A1N(n2137), .Y(n2144)
         );
  AOI2BB2X1 U2260 ( .B0(n2153), .B1(n2152), .A0N(n2153), .A1N(n2151), .Y(n2159) );
  AOI2BB2X1 U2261 ( .B0(n2169), .B1(n2170), .A0N(n2169), .A1N(n2168), .Y(n2181) );
  OAI2BB2XL U2262 ( .B0(n2181), .B1(n2173), .A0N(n2181), .A1N(n2184), .Y(n2185) );
  AOI2BB2X1 U2263 ( .B0(n2178), .B1(n2179), .A0N(n2178), .A1N(n2179), .Y(n2177) );
  OAI21XL U2264 ( .A0(n2175), .A1(n2174), .B0(n2187), .Y(n2176) );
  AOI2BB2X1 U2265 ( .B0(n659), .B1(n2177), .A0N(n2211), .A1N(n2176), .Y(n2229)
         );
  AOI2BB2X1 U2266 ( .B0(curr_photo[0]), .B1(photo_num[0]), .A0N(curr_photo[0]), 
        .A1N(photo_num[0]), .Y(n2217) );
  AOI2BB2X1 U2267 ( .B0(curr_photo[1]), .B1(photo_num[1]), .A0N(curr_photo[1]), 
        .A1N(photo_num[1]), .Y(n2216) );
  OAI21XL U2268 ( .A0(n2234), .A1(N76), .B0(n2239), .Y(n2226) );
  OAI22XL U2269 ( .A0(read_cntr[0]), .A1(n2244), .B0(n277), .B1(n2243), .Y(
        n336) );
endmodule


module DPA ( clk, reset, IM_A, IM_Q, IM_D, IM_WEN, CR_A, CR_Q );
  output [19:0] IM_A;
  input [23:0] IM_Q;
  output [23:0] IM_D;
  output [8:0] CR_A;
  input [12:0] CR_Q;
  input clk, reset;
  output IM_WEN;
  wire   n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, im_d_w_19, im_d_w_18,
         im_d_w_9, im_d_w_8, en_si, en_init_time, en_photo_num,
         en_curr_photo_size, en_so, si_sel, init_time_mux_sel,
         \data_path/si_w[0] , \data_path/si_w[1] , \data_path/si_w[2] ,
         \data_path/si_w[3] , \data_path/si_w[4] , \data_path/si_w[5] ,
         \data_path/si_w[6] , \data_path/si_w[7] , \data_path/si_w[8] ,
         \data_path/si_w[9] , \data_path/si_w[10] , \data_path/si_w[11] ,
         \data_path/si_w[12] , \data_path/si_w[13] , \data_path/si_w[14] ,
         \data_path/si_w[15] , \data_path/si_w[16] , \data_path/si_w[17] ,
         \data_path/si_w[18] , \data_path/si_w[19] , \data_path/si_w[20] ,
         \data_path/si_w[21] , \data_path/si_w[22] , \data_path/si_w[23] , n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n141,
         n144, n145, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         \intadd_0/CI , \intadd_0/SUM[5] , \intadd_0/SUM[4] ,
         \intadd_0/SUM[3] , \intadd_0/SUM[2] , \intadd_0/SUM[1] ,
         \intadd_0/SUM[0] , \intadd_0/CO , \intadd_0/n6 , \intadd_0/n5 ,
         \intadd_0/n4 , \intadd_0/n3 , \intadd_0/n2 , \intadd_0/n1 ,
         \intadd_1/CI , \intadd_1/SUM[5] , \intadd_1/SUM[4] ,
         \intadd_1/SUM[3] , \intadd_1/SUM[2] , \intadd_1/SUM[1] ,
         \intadd_1/SUM[0] , \intadd_1/n6 , \intadd_1/n5 , \intadd_1/n4 ,
         \intadd_1/n3 , \intadd_1/n2 , \intadd_1/n1 , \intadd_2/CI ,
         \intadd_2/SUM[5] , \intadd_2/SUM[4] , \intadd_2/SUM[3] ,
         \intadd_2/SUM[2] , \intadd_2/SUM[1] , \intadd_2/SUM[0] ,
         \intadd_2/CO , \intadd_2/n6 , \intadd_2/n5 , \intadd_2/n4 ,
         \intadd_2/n3 , \intadd_2/n2 , \intadd_2/n1 , n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n431, n433, n435, n437, n439, n440,
         n473, n474, n475, n476, n477, n478, n480, n482, n484, n486, n488,
         n490, n492, n494, n496, n498, n500, n502, n504, n506, n508, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n768;
  wire   [29:28] im_d_w;
  wire   [23:0] curr_time;
  wire   [19:0] fb_addr;
  wire   [1:0] photo_num;
  wire   [19:0] curr_photo_addr;
  wire   [1:0] curr_photo_size;
  wire   [1:0] so_mux_sel;
  wire   [3:0] expand_sel;

  CONT ctrl_logic ( .clk(clk), .reset(reset), .im_wen_n(IM_WEN), .cr_a(CR_A), 
        .curr_time({curr_time[23:10], n477, curr_time[8:0]}), .fb_addr(fb_addr), .photo_num(photo_num), .curr_photo_addr(curr_photo_addr), .curr_photo_size(
        curr_photo_size), .en_si(en_si), .en_init_time(en_init_time), 
        .en_fb_addr(n476), .en_photo_num(en_photo_num), .en_curr_photo_addr(
        n475), .en_curr_photo_size(en_curr_photo_size), .en_so(en_so), 
        .si_sel(si_sel), .init_time_mux_sel(init_time_mux_sel), .so_mux_sel(
        so_mux_sel), .expand_sel(expand_sel), .\im_a[19]_BAR (n769), 
        .\im_a[18]_BAR (n770), .\im_a[17]_BAR (n771), .\im_a[16]_BAR (n772), 
        .\im_a[15]_BAR (n773), .\im_a[14]_BAR (n774), .\im_a[13]_BAR (n775), 
        .\im_a[12]_BAR (n776), .\im_a[11]_BAR (n777), .\im_a[10]_BAR (n778), 
        .\im_a[9]_BAR (n779), .\im_a[8]_BAR (n780), .\im_a[7]_BAR (n781), 
        .\im_a[6]_BAR (n782), .\im_a[5]_BAR (n783), .\im_a[4]_BAR (n784), 
        .\im_a[3]_BAR (n785), .\im_a[2]_BAR (n786), .\im_a[1]_BAR (n787), 
        .\im_a[0]_BAR (n788) );
  ADDFXL \intadd_0/U3  ( .A(n790), .B(\data_path/si_w[22] ), .CI(\intadd_0/n3 ), .CO(\intadd_0/n2 ), .S(\intadd_0/SUM[4] ) );
  DFFSX1 \data_path/init_time_reg/q_reg[1]  ( .D(n145), .CK(clk), .SN(n439), 
        .Q(n515), .QN(curr_time[1]) );
  CLKBUFX3 \intadd_2/U1  ( .A(\intadd_2/n1 ), .Y(\intadd_2/CO ) );
  CLKBUFX3 \intadd_0/U1  ( .A(\intadd_0/n1 ), .Y(\intadd_0/CO ) );
  ADDFXL \intadd_0/U5  ( .A(n792), .B(\data_path/si_w[20] ), .CI(\intadd_0/n5 ), .CO(\intadd_0/n4 ), .S(\intadd_0/SUM[2] ) );
  ADDFXL \intadd_0/U2  ( .A(n789), .B(\data_path/si_w[23] ), .CI(\intadd_0/n2 ), .CO(\intadd_0/n1 ), .S(\intadd_0/SUM[5] ) );
  ADDFXL \intadd_1/U7  ( .A(IM_D[10]), .B(\data_path/si_w[10] ), .CI(
        \intadd_1/CI ), .CO(\intadd_1/n6 ), .S(\intadd_1/SUM[0] ) );
  ADDFXL \intadd_1/U3  ( .A(IM_D[14]), .B(\data_path/si_w[14] ), .CI(
        \intadd_1/n3 ), .CO(\intadd_1/n2 ), .S(\intadd_1/SUM[4] ) );
  ADDFXL \intadd_1/U2  ( .A(IM_D[15]), .B(\data_path/si_w[15] ), .CI(
        \intadd_1/n2 ), .CO(\intadd_1/n1 ), .S(\intadd_1/SUM[5] ) );
  ADDFXL \intadd_2/U7  ( .A(IM_D[2]), .B(\data_path/si_w[2] ), .CI(
        \intadd_2/CI ), .CO(\intadd_2/n6 ), .S(\intadd_2/SUM[0] ) );
  ADDFXL \intadd_2/U3  ( .A(IM_D[6]), .B(\data_path/si_w[6] ), .CI(
        \intadd_2/n3 ), .CO(\intadd_2/n2 ), .S(\intadd_2/SUM[4] ) );
  ADDFXL \intadd_2/U2  ( .A(IM_D[7]), .B(\data_path/si_w[7] ), .CI(
        \intadd_2/n2 ), .CO(\intadd_2/n1 ), .S(\intadd_2/SUM[5] ) );
  ADDFXL \intadd_0/U7  ( .A(IM_D[18]), .B(\data_path/si_w[18] ), .CI(
        \intadd_0/CI ), .CO(\intadd_0/n6 ), .S(\intadd_0/SUM[0] ) );
  ADDFXL \intadd_0/U4  ( .A(n791), .B(\data_path/si_w[21] ), .CI(\intadd_0/n4 ), .CO(\intadd_0/n3 ), .S(\intadd_0/SUM[3] ) );
  ADDFXL \intadd_0/U6  ( .A(n793), .B(\data_path/si_w[19] ), .CI(\intadd_0/n6 ), .CO(\intadd_0/n5 ), .S(\intadd_0/SUM[1] ) );
  ADDFXL \intadd_1/U6  ( .A(IM_D[11]), .B(\data_path/si_w[11] ), .CI(
        \intadd_1/n6 ), .CO(\intadd_1/n5 ), .S(\intadd_1/SUM[1] ) );
  ADDFXL \intadd_2/U6  ( .A(IM_D[3]), .B(\data_path/si_w[3] ), .CI(
        \intadd_2/n6 ), .CO(\intadd_2/n5 ), .S(\intadd_2/SUM[1] ) );
  DFFSX2 \data_path/si_reg/q_reg[8]  ( .D(n312), .CK(clk), .SN(n22), .Q(n520), 
        .QN(\data_path/si_w[8] ) );
  ADDFXL \intadd_1/U5  ( .A(IM_D[12]), .B(\data_path/si_w[12] ), .CI(
        \intadd_1/n5 ), .CO(\intadd_1/n4 ), .S(\intadd_1/SUM[2] ) );
  ADDFXL \intadd_1/U4  ( .A(IM_D[13]), .B(\data_path/si_w[13] ), .CI(
        \intadd_1/n4 ), .CO(\intadd_1/n3 ), .S(\intadd_1/SUM[3] ) );
  ADDFXL \intadd_2/U5  ( .A(IM_D[4]), .B(\data_path/si_w[4] ), .CI(
        \intadd_2/n5 ), .CO(\intadd_2/n4 ), .S(\intadd_2/SUM[2] ) );
  ADDFXL \intadd_2/U4  ( .A(IM_D[5]), .B(\data_path/si_w[5] ), .CI(
        \intadd_2/n4 ), .CO(\intadd_2/n3 ), .S(\intadd_2/SUM[3] ) );
  DFFSX2 \data_path/si_reg/q_reg[4]  ( .D(n313), .CK(clk), .SN(n22), .QN(
        \data_path/si_w[4] ) );
  DFFSX2 \data_path/si_reg/q_reg[2]  ( .D(n314), .CK(clk), .SN(n439), .QN(
        \data_path/si_w[2] ) );
  DFFSX2 \data_path/si_reg/q_reg[1]  ( .D(n315), .CK(clk), .SN(n440), .Q(n745), 
        .QN(\data_path/si_w[1] ) );
  DFFSX2 \data_path/init_time_reg/q_reg[2]  ( .D(n144), .CK(clk), .SN(n22), 
        .QN(curr_time[2]) );
  DFFSX2 \data_path/init_time_reg/q_reg[4]  ( .D(n141), .CK(clk), .SN(n439), 
        .QN(curr_time[4]) );
  DFFRX1 \data_path/si_reg/q_reg[22]  ( .D(n370), .CK(clk), .RN(n440), .Q(
        \data_path/si_w[22] ) );
  DFFRX1 \data_path/si_reg/q_reg[21]  ( .D(n371), .CK(clk), .RN(n439), .Q(
        \data_path/si_w[21] ) );
  DFFRX1 \data_path/si_reg/q_reg[20]  ( .D(n372), .CK(clk), .RN(n22), .Q(
        \data_path/si_w[20] ) );
  DFFRX1 \data_path/photo_num_reg/q_reg[0]  ( .D(n367), .CK(clk), .RN(n440), 
        .Q(photo_num[0]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[18]  ( .D(n377), .CK(clk), .RN(n439), 
        .Q(fb_addr[18]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[13]  ( .D(n389), .CK(clk), .RN(n22), .Q(
        fb_addr[13]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[18]  ( .D(n376), .CK(clk), .RN(
        n440), .Q(curr_photo_addr[18]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[13]  ( .D(n388), .CK(clk), .RN(
        n439), .Q(curr_photo_addr[13]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[15]  ( .D(n383), .CK(clk), .RN(n22), .Q(
        fb_addr[15]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[14]  ( .D(n386), .CK(clk), .RN(n440), 
        .Q(fb_addr[14]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[9]  ( .D(n401), .CK(clk), .RN(n439), .Q(
        fb_addr[9]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[8]  ( .D(n14), .CK(clk), .RN(n22), .Q(
        fb_addr[8]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[7]  ( .D(n404), .CK(clk), .RN(n440), .Q(
        fb_addr[7]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[3]  ( .D(n413), .CK(clk), .RN(n439), .Q(
        fb_addr[3]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[0]  ( .D(n416), .CK(clk), .RN(n22), .Q(
        fb_addr[0]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[19]  ( .D(n374), .CK(clk), .RN(n440), 
        .Q(fb_addr[19]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[12]  ( .D(n392), .CK(clk), .RN(n439), 
        .Q(fb_addr[12]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[10]  ( .D(n398), .CK(clk), .RN(n22), .Q(
        fb_addr[10]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[6]  ( .D(n407), .CK(clk), .RN(n440), .Q(
        fb_addr[6]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[5]  ( .D(n410), .CK(clk), .RN(n439), .Q(
        fb_addr[5]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[17]  ( .D(n380), .CK(clk), .RN(n22), .Q(
        fb_addr[17]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[11]  ( .D(n395), .CK(clk), .RN(n440), 
        .Q(fb_addr[11]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[1]  ( .D(n20), .CK(clk), .RN(n439), .Q(
        fb_addr[1]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[9]  ( .D(n400), .CK(clk), .RN(
        n22), .Q(curr_photo_addr[9]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[8]  ( .D(n13), .CK(clk), .RN(
        n440), .Q(curr_photo_addr[8]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[7]  ( .D(n403), .CK(clk), .RN(
        n439), .Q(curr_photo_addr[7]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[3]  ( .D(n412), .CK(clk), .RN(
        n22), .Q(curr_photo_addr[3]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[15]  ( .D(n382), .CK(clk), .RN(
        n440), .Q(curr_photo_addr[15]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[14]  ( .D(n385), .CK(clk), .RN(
        n439), .Q(curr_photo_addr[14]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[0]  ( .D(n415), .CK(clk), .RN(
        n22), .Q(curr_photo_addr[0]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[19]  ( .D(n373), .CK(clk), .RN(
        n440), .Q(curr_photo_addr[19]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[12]  ( .D(n391), .CK(clk), .RN(
        n439), .Q(curr_photo_addr[12]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[10]  ( .D(n397), .CK(clk), .RN(
        n22), .Q(curr_photo_addr[10]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[6]  ( .D(n406), .CK(clk), .RN(
        n440), .Q(curr_photo_addr[6]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[5]  ( .D(n409), .CK(clk), .RN(
        n439), .Q(curr_photo_addr[5]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[17]  ( .D(n379), .CK(clk), .RN(
        n22), .Q(curr_photo_addr[17]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[11]  ( .D(n394), .CK(clk), .RN(
        n440), .Q(curr_photo_addr[11]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[1]  ( .D(n19), .CK(clk), .RN(
        n439), .Q(curr_photo_addr[1]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[16]  ( .D(n12), .CK(clk), .RN(n22), .Q(
        fb_addr[16]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[16]  ( .D(n11), .CK(clk), .RN(
        n440), .Q(curr_photo_addr[16]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[4]  ( .D(n16), .CK(clk), .RN(n439), .Q(
        fb_addr[4]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[2]  ( .D(n18), .CK(clk), .RN(n22), .Q(
        fb_addr[2]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[4]  ( .D(n15), .CK(clk), .RN(
        n440), .Q(curr_photo_addr[4]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[2]  ( .D(n17), .CK(clk), .RN(
        n439), .Q(curr_photo_addr[2]) );
  DFFRX1 \data_path/init_time_reg/q_reg[21]  ( .D(n318), .CK(clk), .RN(n22), 
        .Q(curr_time[21]) );
  DFFRX1 \data_path/init_time_reg/q_reg[5]  ( .D(n334), .CK(clk), .RN(n440), 
        .Q(curr_time[5]) );
  DFFRX1 \data_path/init_time_reg/q_reg[8]  ( .D(n331), .CK(clk), .RN(n439), 
        .Q(curr_time[8]) );
  DFFRX1 \data_path/so_reg/q_reg[29]  ( .D(n337), .CK(clk), .RN(n22), .Q(
        im_d_w[29]) );
  DFFRX1 \data_path/so_reg/q_reg[19]  ( .D(n347), .CK(clk), .RN(n440), .Q(
        im_d_w_19) );
  DFFRX1 \data_path/so_reg/q_reg[18]  ( .D(n348), .CK(clk), .RN(n439), .Q(
        im_d_w_18) );
  DFFRX1 \data_path/so_reg/q_reg[9]  ( .D(n357), .CK(clk), .RN(n22), .Q(
        im_d_w_9) );
  DFFRX1 \data_path/so_reg/q_reg[0]  ( .D(n366), .CK(clk), .RN(n440), .QN(n508) );
  DFFRX1 \data_path/so_reg/q_reg[15]  ( .D(n351), .CK(clk), .RN(n439), .QN(
        n504) );
  DFFRX1 \data_path/so_reg/q_reg[14]  ( .D(n352), .CK(clk), .RN(n22), .QN(n498) );
  DFFRX1 \data_path/so_reg/q_reg[5]  ( .D(n361), .CK(clk), .RN(n440), .QN(n506) );
  DFFRX1 \data_path/so_reg/q_reg[4]  ( .D(n362), .CK(clk), .RN(n439), .QN(n500) );
  DFFRX1 \data_path/so_reg/q_reg[3]  ( .D(n363), .CK(clk), .RN(n22), .QN(n502)
         );
  DFFRX1 \data_path/so_reg/q_reg[17]  ( .D(n349), .CK(clk), .RN(n440), .QN(
        n490) );
  DFFRX1 \data_path/so_reg/q_reg[16]  ( .D(n350), .CK(clk), .RN(n439), .QN(
        n488) );
  DFFRX1 \data_path/so_reg/q_reg[7]  ( .D(n359), .CK(clk), .RN(n22), .QN(n492)
         );
  DFFRX1 \data_path/so_reg/q_reg[6]  ( .D(n360), .CK(clk), .RN(n440), .QN(n494) );
  DFFRX1 \data_path/so_reg/q_reg[22]  ( .D(n344), .CK(clk), .RN(n439), .QN(
        n486) );
  DFFRX1 \data_path/so_reg/q_reg[2]  ( .D(n364), .CK(clk), .RN(n22), .QN(n496)
         );
  DFFRX1 \data_path/si_reg/q_reg[9]  ( .D(n402), .CK(clk), .RN(n440), .Q(
        \data_path/si_w[9] ), .QN(n527) );
  DFFRX1 \data_path/init_time_reg/q_reg[9]  ( .D(n330), .CK(clk), .RN(n440), 
        .Q(curr_time[9]), .QN(n539) );
  DFFRX1 \data_path/so_reg/q_reg[11]  ( .D(n355), .CK(clk), .RN(n440), .QN(
        n480) );
  DFFSRX1 \data_path/si_reg/q_reg[23]  ( .D(n369), .CK(clk), .SN(1'b1), .RN(
        n439), .Q(\data_path/si_w[23] ), .QN(n526) );
  DFFSRX1 \data_path/si_reg/q_reg[19]  ( .D(n375), .CK(clk), .SN(1'b1), .RN(
        n22), .Q(\data_path/si_w[19] ), .QN(n538) );
  DFFSRX1 \data_path/si_reg/q_reg[18]  ( .D(n378), .CK(clk), .SN(1'b1), .RN(
        n440), .Q(\data_path/si_w[18] ), .QN(n535) );
  DFFSRX1 \data_path/si_reg/q_reg[17]  ( .D(n381), .CK(clk), .SN(1'b1), .RN(
        n439), .Q(\data_path/si_w[17] ), .QN(n528) );
  DFFSRX1 \data_path/si_reg/q_reg[15]  ( .D(n384), .CK(clk), .SN(1'b1), .RN(
        n22), .Q(\data_path/si_w[15] ), .QN(n542) );
  DFFSRX1 \data_path/si_reg/q_reg[14]  ( .D(n387), .CK(clk), .SN(1'b1), .RN(
        n440), .Q(\data_path/si_w[14] ), .QN(n541) );
  DFFSRX1 \data_path/si_reg/q_reg[13]  ( .D(n390), .CK(clk), .SN(1'b1), .RN(
        n439), .Q(\data_path/si_w[13] ), .QN(n523) );
  DFFSRX1 \data_path/si_reg/q_reg[12]  ( .D(n393), .CK(clk), .SN(1'b1), .RN(
        n22), .Q(\data_path/si_w[12] ), .QN(n533) );
  DFFSRX1 \data_path/si_reg/q_reg[11]  ( .D(n396), .CK(clk), .SN(1'b1), .RN(
        n440), .Q(\data_path/si_w[11] ), .QN(n517) );
  DFFSRX1 \data_path/si_reg/q_reg[10]  ( .D(n399), .CK(clk), .SN(1'b1), .RN(
        n439), .Q(\data_path/si_w[10] ), .QN(n514) );
  DFFSRX1 \data_path/si_reg/q_reg[6]  ( .D(n408), .CK(clk), .SN(1'b1), .RN(n22), .Q(\data_path/si_w[6] ), .QN(n534) );
  DFFSRX1 \data_path/si_reg/q_reg[5]  ( .D(n411), .CK(clk), .SN(1'b1), .RN(
        n440), .Q(\data_path/si_w[5] ), .QN(n524) );
  DFFSRX1 \data_path/photo_num_reg/q_reg[1]  ( .D(n21), .CK(clk), .SN(1'b1), 
        .RN(n439), .Q(photo_num[1]), .QN(n10) );
  DFFSRX1 \data_path/init_time_reg/q_reg[16]  ( .D(n323), .CK(clk), .SN(1'b1), 
        .RN(n22), .Q(curr_time[16]), .QN(n518) );
  DFFSRX1 \data_path/curr_photo_size_reg/q_reg[1]  ( .D(n23), .CK(clk), .SN(
        1'b1), .RN(n440), .Q(curr_photo_size[1]), .QN(n547) );
  DFFSRX1 \data_path/curr_photo_size_reg/q_reg[0]  ( .D(n368), .CK(clk), .SN(
        1'b1), .RN(n439), .Q(curr_photo_size[0]), .QN(n525) );
  DFFSRX1 \data_path/init_time_reg/q_reg[3]  ( .D(n335), .CK(clk), .SN(1'b1), 
        .RN(n22), .Q(curr_time[3]), .QN(n540) );
  DFFSRX1 \data_path/init_time_reg/q_reg[0]  ( .D(n336), .CK(clk), .SN(1'b1), 
        .RN(n440), .Q(curr_time[0]), .QN(n529) );
  DFFSRX1 \data_path/init_time_reg/q_reg[11]  ( .D(n328), .CK(clk), .SN(1'b1), 
        .RN(n439), .Q(curr_time[11]), .QN(n516) );
  DFFSRX1 \data_path/init_time_reg/q_reg[13]  ( .D(n326), .CK(clk), .SN(1'b1), 
        .RN(n22), .Q(curr_time[13]), .QN(n545) );
  DFFSRX1 \data_path/init_time_reg/q_reg[23]  ( .D(n316), .CK(clk), .SN(1'b1), 
        .RN(n440), .Q(curr_time[23]), .QN(n519) );
  DFFSRX1 \data_path/init_time_reg/q_reg[19]  ( .D(n320), .CK(clk), .SN(1'b1), 
        .RN(n439), .Q(curr_time[19]), .QN(n546) );
  DFFSRX1 \data_path/init_time_reg/q_reg[10]  ( .D(n329), .CK(clk), .SN(1'b1), 
        .RN(n22), .Q(curr_time[10]), .QN(n521) );
  DFFSRX1 \data_path/so_reg/q_reg[28]  ( .D(n338), .CK(clk), .SN(1'b1), .RN(
        n440), .Q(im_d_w[28]), .QN(n544) );
  DFFSRX1 \data_path/so_reg/q_reg[8]  ( .D(n358), .CK(clk), .SN(1'b1), .RN(
        n439), .Q(im_d_w_8), .QN(n543) );
  DFFSRX1 \data_path/so_reg/q_reg[25]  ( .D(n341), .CK(clk), .SN(1'b1), .RN(
        n22), .Q(n791), .QN(n435) );
  DFFSRX1 \data_path/so_reg/q_reg[24]  ( .D(n342), .CK(clk), .SN(1'b1), .RN(
        n440), .Q(n792), .QN(n437) );
  DFFSRX1 \data_path/so_reg/q_reg[21]  ( .D(n345), .CK(clk), .SN(1'b1), .RN(
        n439), .QN(n482) );
  DFFSRX1 \data_path/so_reg/q_reg[1]  ( .D(n365), .CK(clk), .SN(1'b1), .RN(n22), .QN(n484) );
  DFFSRX1 \data_path/so_reg/q_reg[23]  ( .D(n343), .CK(clk), .SN(1'b1), .RN(
        n440), .Q(n793), .QN(n429) );
  DFFSRX1 \data_path/so_reg/q_reg[27]  ( .D(n339), .CK(clk), .SN(1'b1), .RN(
        n439), .Q(n789), .QN(n433) );
  DFFSRX1 \data_path/so_reg/q_reg[26]  ( .D(n340), .CK(clk), .SN(1'b1), .RN(
        n440), .Q(n790), .QN(n431) );
  DFFRX2 \data_path/si_reg/q_reg[16]  ( .D(n418), .CK(clk), .RN(n22), .Q(
        \data_path/si_w[16] ) );
  DFFRX2 \data_path/init_time_reg/q_reg[15]  ( .D(n324), .CK(clk), .RN(n439), 
        .Q(curr_time[15]) );
  DFFRX2 \data_path/init_time_reg/q_reg[14]  ( .D(n325), .CK(clk), .RN(n439), 
        .Q(curr_time[14]) );
  DFFRX2 \data_path/init_time_reg/q_reg[7]  ( .D(n332), .CK(clk), .RN(n439), 
        .Q(curr_time[7]) );
  DFFRX2 \data_path/init_time_reg/q_reg[6]  ( .D(n333), .CK(clk), .RN(n22), 
        .Q(curr_time[6]) );
  DFFRX2 \data_path/init_time_reg/q_reg[22]  ( .D(n317), .CK(clk), .RN(n22), 
        .Q(curr_time[22]) );
  DFFRX2 \data_path/init_time_reg/q_reg[20]  ( .D(n319), .CK(clk), .RN(n439), 
        .Q(curr_time[20]) );
  DFFRX2 \data_path/si_reg/q_reg[0]  ( .D(n417), .CK(clk), .RN(n440), .Q(
        \data_path/si_w[0] ), .QN(n531) );
  DFFRX2 \data_path/init_time_reg/q_reg[17]  ( .D(n322), .CK(clk), .RN(n22), 
        .Q(curr_time[17]), .QN(n532) );
  DFFRX2 \data_path/init_time_reg/q_reg[18]  ( .D(n321), .CK(clk), .RN(n439), 
        .Q(curr_time[18]), .QN(n522) );
  DFFRX2 \data_path/init_time_reg/q_reg[12]  ( .D(n327), .CK(clk), .RN(n22), 
        .Q(curr_time[12]), .QN(n530) );
  DFFRX2 \data_path/si_reg/q_reg[3]  ( .D(n414), .CK(clk), .RN(n22), .Q(
        \data_path/si_w[3] ), .QN(n537) );
  DFFRX2 \data_path/si_reg/q_reg[7]  ( .D(n405), .CK(clk), .RN(n439), .Q(
        \data_path/si_w[7] ), .QN(n536) );
  DFFRX1 \data_path/so_reg/q_reg[20]  ( .D(n346), .CK(clk), .RN(n439), .Q(n794) );
  DFFRX1 \data_path/so_reg/q_reg[10]  ( .D(n356), .CK(clk), .RN(n22), .Q(n797)
         );
  DFFRX1 \data_path/so_reg/q_reg[13]  ( .D(n353), .CK(clk), .RN(n439), .Q(n795) );
  DFFRX1 \data_path/so_reg/q_reg[12]  ( .D(n354), .CK(clk), .RN(n22), .Q(n796)
         );
  BUFX4 U435 ( .A(n743), .Y(n549) );
  CLKBUFX3 U436 ( .A(n744), .Y(n550) );
  NOR4X1 U437 ( .A(\data_path/si_w[16] ), .B(\data_path/si_w[17] ), .C(
        \data_path/si_w[18] ), .D(\data_path/si_w[19] ), .Y(n421) );
  NOR4X1 U438 ( .A(\data_path/si_w[1] ), .B(\data_path/si_w[2] ), .C(
        \data_path/si_w[15] ), .D(\data_path/si_w[23] ), .Y(n422) );
  NOR4X1 U439 ( .A(\data_path/si_w[20] ), .B(\data_path/si_w[14] ), .C(
        \data_path/si_w[21] ), .D(\data_path/si_w[22] ), .Y(n423) );
  AND4X1 U440 ( .A(n523), .B(n520), .C(n533), .D(en_curr_photo_size), .Y(n424)
         );
  AND4X1 U441 ( .A(n421), .B(n422), .C(n423), .D(n424), .Y(n558) );
  CLKINVX1 U442 ( .A(n475), .Y(n551) );
  OAI2BB1X1 U443 ( .A0N(IM_D[8]), .A1N(\data_path/si_w[8] ), .B0(n527), .Y(
        n608) );
  CLKINVX1 U444 ( .A(n476), .Y(n552) );
  NAND2X1 U445 ( .A(n543), .B(\intadd_2/CO ), .Y(n425) );
  AOI2BB1X1 U446 ( .A0N(\intadd_2/CO ), .A1N(n707), .B0(n740), .Y(n426) );
  OAI22XL U447 ( .A0(n741), .A1(n425), .B0(n426), .B1(n543), .Y(n358) );
  NAND3BX1 U448 ( .AN(n527), .B(IM_D[8]), .C(\data_path/si_w[8] ), .Y(n607) );
  AOI2BB1X1 U449 ( .A0N(\intadd_0/CO ), .A1N(n707), .B0(n740), .Y(n427) );
  NAND2X1 U450 ( .A(n544), .B(\intadd_0/CO ), .Y(n428) );
  OAI22XL U451 ( .A0(n741), .A1(n428), .B0(n427), .B1(n544), .Y(n338) );
  AOI211X1 U452 ( .A0(curr_time[13]), .A1(n683), .B0(curr_time[15]), .C0(
        curr_time[14]), .Y(n690) );
  INVX16 U453 ( .A(n429), .Y(IM_D[19]) );
  INVX16 U454 ( .A(n431), .Y(IM_D[22]) );
  INVX16 U455 ( .A(n433), .Y(IM_D[23]) );
  INVX16 U456 ( .A(n435), .Y(IM_D[21]) );
  INVX16 U457 ( .A(n437), .Y(IM_D[20]) );
  INVX8 U458 ( .A(reset), .Y(n439) );
  INVX6 U459 ( .A(reset), .Y(n440) );
  INVX8 U460 ( .A(reset), .Y(n22) );
  NOR2X1 U493 ( .A(n671), .B(n673), .Y(n679) );
  INVX6 U494 ( .A(n551), .Y(n473) );
  INVX6 U495 ( .A(n552), .Y(n474) );
  INVX6 U496 ( .A(en_so), .Y(n740) );
  INVX3 U497 ( .A(en_si), .Y(n744) );
  NOR2X1 U498 ( .A(si_sel), .B(n550), .Y(n743) );
  BUFX2 U499 ( .A(curr_time[9]), .Y(n477) );
  NOR2X1 U500 ( .A(n540), .B(n671), .Y(n674) );
  NAND2X1 U501 ( .A(curr_time[2]), .B(n668), .Y(n671) );
  CLKINVX1 U502 ( .A(n663), .Y(n673) );
  NOR2X1 U503 ( .A(n684), .B(n677), .Y(n663) );
  NAND2BX1 U504 ( .AN(n737), .B(n686), .Y(n706) );
  NAND2X1 U505 ( .A(n688), .B(n690), .Y(n686) );
  NOR2X1 U506 ( .A(n518), .B(n699), .Y(n694) );
  NAND2X1 U507 ( .A(en_init_time), .B(n692), .Y(n699) );
  INVX3 U508 ( .A(n741), .Y(n658) );
  CLKINVX1 U509 ( .A(n692), .Y(n700) );
  AOI211X1 U510 ( .A0(n701), .A1(curr_time[20]), .B0(n690), .C0(n689), .Y(n692) );
  AOI211X1 U511 ( .A0(n661), .A1(curr_time[5]), .B0(curr_time[6]), .C0(
        curr_time[7]), .Y(n682) );
  NOR2X1 U512 ( .A(curr_time[8]), .B(n728), .Y(n713) );
  OAI221XL U513 ( .A0(expand_sel[0]), .A1(\data_path/si_w[8] ), .B0(n570), 
        .B1(\data_path/si_w[7] ), .C0(n573), .Y(n569) );
  CLKINVX1 U514 ( .A(n548), .Y(n629) );
  BUFX4 U515 ( .A(n655), .Y(n548) );
  NOR2X1 U516 ( .A(curr_time[2]), .B(n668), .Y(n666) );
  AOI211X1 U517 ( .A0(curr_time[2]), .A1(n668), .B0(n684), .C0(n677), .Y(n669)
         );
  NOR2X2 U518 ( .A(n515), .B(n529), .Y(n668) );
  CLKINVX1 U519 ( .A(expand_sel[1]), .Y(n573) );
  INVX3 U520 ( .A(n660), .Y(n647) );
  NAND3X2 U521 ( .A(so_mux_sel[0]), .B(so_mux_sel[1]), .C(en_so), .Y(n660) );
  INVX16 U522 ( .A(n788), .Y(IM_A[0]) );
  INVX16 U523 ( .A(n787), .Y(IM_A[1]) );
  INVX16 U524 ( .A(n786), .Y(IM_A[2]) );
  INVX16 U525 ( .A(n785), .Y(IM_A[3]) );
  INVX16 U526 ( .A(n784), .Y(IM_A[4]) );
  INVX16 U527 ( .A(n783), .Y(IM_A[5]) );
  INVX16 U528 ( .A(n782), .Y(IM_A[6]) );
  INVX16 U529 ( .A(n781), .Y(IM_A[7]) );
  INVX16 U530 ( .A(n780), .Y(IM_A[8]) );
  INVX16 U531 ( .A(n779), .Y(IM_A[9]) );
  INVX16 U532 ( .A(n778), .Y(IM_A[10]) );
  INVX16 U533 ( .A(n777), .Y(IM_A[11]) );
  INVX16 U534 ( .A(n776), .Y(IM_A[12]) );
  INVX16 U535 ( .A(n775), .Y(IM_A[13]) );
  INVX16 U536 ( .A(n774), .Y(IM_A[14]) );
  INVX16 U537 ( .A(n773), .Y(IM_A[15]) );
  INVX16 U538 ( .A(n772), .Y(IM_A[16]) );
  INVX16 U539 ( .A(n771), .Y(IM_A[17]) );
  INVX16 U540 ( .A(n770), .Y(IM_A[18]) );
  CLKINVX1 U541 ( .A(n768), .Y(n478) );
  INVX16 U542 ( .A(n478), .Y(IM_A[19]) );
  INVX16 U543 ( .A(n480), .Y(IM_D[9]) );
  INVX16 U544 ( .A(n482), .Y(IM_D[17]) );
  INVX16 U545 ( .A(n484), .Y(IM_D[1]) );
  INVX16 U546 ( .A(n486), .Y(IM_D[18]) );
  INVX16 U547 ( .A(n488), .Y(IM_D[14]) );
  INVX16 U548 ( .A(n490), .Y(IM_D[15]) );
  INVX16 U549 ( .A(n492), .Y(IM_D[7]) );
  INVX16 U550 ( .A(n494), .Y(IM_D[6]) );
  INVX16 U551 ( .A(n496), .Y(IM_D[2]) );
  INVX16 U552 ( .A(n498), .Y(IM_D[12]) );
  INVX16 U553 ( .A(n500), .Y(IM_D[4]) );
  INVX16 U554 ( .A(n502), .Y(IM_D[3]) );
  INVX16 U555 ( .A(n504), .Y(IM_D[13]) );
  INVX16 U556 ( .A(n506), .Y(IM_D[5]) );
  INVX16 U557 ( .A(n508), .Y(IM_D[0]) );
  NOR2X1 U558 ( .A(n521), .B(n722), .Y(n723) );
  OAI21X1 U559 ( .A0(\intadd_1/n1 ), .A1(im_d_w_18), .B0(n625), .Y(n739) );
  NAND2X1 U560 ( .A(\intadd_1/n1 ), .B(im_d_w_18), .Y(n625) );
  NOR2X1 U561 ( .A(\data_path/si_w[4] ), .B(n556), .Y(n559) );
  NOR2X1 U562 ( .A(n713), .B(n737), .Y(n717) );
  NAND2X2 U563 ( .A(en_init_time), .B(n677), .Y(n737) );
  NOR2BX1 U564 ( .AN(init_time_mux_sel), .B(n682), .Y(n688) );
  NAND2X1 U565 ( .A(n682), .B(init_time_mux_sel), .Y(n677) );
  CLKINVX1 U566 ( .A(n724), .Y(n728) );
  NAND2X1 U567 ( .A(n724), .B(n723), .Y(n733) );
  NOR2X1 U568 ( .A(n686), .B(n684), .Y(n724) );
  NAND3XL U569 ( .A(\data_path/si_w[0] ), .B(\data_path/si_w[1] ), .C(IM_D[0]), 
        .Y(n582) );
  NOR2BX1 U570 ( .AN(n701), .B(n699), .Y(n703) );
  NOR3X2 U571 ( .A(n532), .B(n518), .C(n522), .Y(n701) );
  OAI21X1 U572 ( .A0(n701), .A1(n700), .B0(n735), .Y(n704) );
  OAI21X1 U573 ( .A0(curr_time[16]), .A1(n700), .B0(n735), .Y(n695) );
  CLKINVX1 U574 ( .A(n706), .Y(n735) );
  INVX3 U575 ( .A(n648), .Y(n657) );
  OAI211X4 U576 ( .A0(expand_sel[3]), .A1(n580), .B0(n579), .C0(n578), .Y(n648) );
  NOR2X4 U577 ( .A(init_time_mux_sel), .B(n684), .Y(n738) );
  INVX3 U578 ( .A(en_init_time), .Y(n684) );
  CLKINVX1 U579 ( .A(n707), .Y(n554) );
  NAND2BX2 U580 ( .AN(so_mux_sel[1]), .B(so_mux_sel[0]), .Y(n707) );
  CLKINVX1 U581 ( .A(expand_sel[0]), .Y(n570) );
  NOR2X1 U582 ( .A(expand_sel[1]), .B(expand_sel[0]), .Y(n577) );
  BUFX16 U583 ( .A(n796), .Y(IM_D[10]) );
  BUFX16 U584 ( .A(n795), .Y(IM_D[11]) );
  AOI22XL U585 ( .A0(\data_path/si_w[20] ), .A1(n548), .B0(n792), .B1(n740), 
        .Y(n646) );
  AOI22XL U586 ( .A0(n791), .A1(n740), .B0(\data_path/si_w[21] ), .B1(n548), 
        .Y(n650) );
  BUFX16 U587 ( .A(n794), .Y(IM_D[16]) );
  AOI22XL U588 ( .A0(\data_path/si_w[16] ), .A1(n631), .B0(IM_D[16]), .B1(n630), .Y(n632) );
  NAND2XL U589 ( .A(\data_path/si_w[16] ), .B(IM_D[16]), .Y(n628) );
  NAND3XL U590 ( .A(\data_path/si_w[17] ), .B(\data_path/si_w[16] ), .C(
        IM_D[16]), .Y(n633) );
  BUFX16 U591 ( .A(n797), .Y(IM_D[8]) );
  AOI22XL U592 ( .A0(\data_path/si_w[8] ), .A1(n605), .B0(IM_D[8]), .B1(n604), 
        .Y(n606) );
  INVXL U593 ( .A(n732), .Y(n393) );
  INVXL U594 ( .A(n555), .Y(n417) );
  INVXL U595 ( .A(n721), .Y(n399) );
  INVXL U596 ( .A(n726), .Y(n396) );
  INVXL U597 ( .A(n712), .Y(n405) );
  INVXL U598 ( .A(n710), .Y(n411) );
  INVXL U599 ( .A(n711), .Y(n408) );
  INVXL U600 ( .A(n709), .Y(n414) );
  INVXL U601 ( .A(n716), .Y(n402) );
  INVXL U602 ( .A(en_photo_num), .Y(n747) );
  OAI211XL U603 ( .A0(en_curr_photo_size), .A1(n525), .B0(n561), .C0(n748), 
        .Y(n368) );
  NAND4XL U604 ( .A(\data_path/si_w[7] ), .B(n559), .C(n558), .D(n557), .Y(
        n561) );
  NAND4XL U605 ( .A(n560), .B(n559), .C(n558), .D(n536), .Y(n748) );
  INVXL U606 ( .A(n666), .Y(n667) );
  INVXL U607 ( .A(n681), .Y(n334) );
  INVXL U608 ( .A(n678), .Y(n680) );
  AOI211XL U609 ( .A0(curr_time[4]), .A1(n684), .B0(n676), .C0(n675), .Y(n141)
         );
  NOR2BXL U610 ( .AN(\data_path/si_w[4] ), .B(n736), .Y(n675) );
  AOI211XL U611 ( .A0(curr_time[4]), .A1(n674), .B0(n673), .C0(n672), .Y(n676)
         );
  NOR2XL U612 ( .A(curr_time[4]), .B(n674), .Y(n672) );
  OAI32XL U613 ( .A0(n540), .A1(n669), .A2(n684), .B0(n679), .B1(curr_time[3]), 
        .Y(n670) );
  NAND2XL U614 ( .A(curr_time[12]), .B(curr_time[11]), .Y(n734) );
  AOI21XL U615 ( .A0(curr_time[8]), .A1(n737), .B0(n713), .Y(n685) );
  NOR2XL U616 ( .A(n665), .B(n664), .Y(n145) );
  AOI211XL U617 ( .A0(n515), .A1(n529), .B0(n668), .C0(n673), .Y(n665) );
  OAI211XL U618 ( .A0(n736), .A1(n535), .B0(n698), .C0(n697), .Y(n321) );
  NOR2XL U619 ( .A(n700), .B(curr_time[17]), .Y(n696) );
  NAND3XL U620 ( .A(curr_time[17]), .B(n694), .C(n522), .Y(n698) );
  INVXL U621 ( .A(n705), .Y(n319) );
  AOI22XL U622 ( .A0(curr_time[12]), .A1(n729), .B0(n738), .B1(
        \data_path/si_w[12] ), .Y(n730) );
  NAND3XL U623 ( .A(n688), .B(n687), .C(n519), .Y(n689) );
  AOI211XL U624 ( .A0(curr_time[20]), .A1(curr_time[19]), .B0(curr_time[21]), 
        .C0(curr_time[22]), .Y(n687) );
  CLKINVX2 U625 ( .A(n738), .Y(n736) );
  AOI22XL U626 ( .A0(curr_time[10]), .A1(n718), .B0(\data_path/si_w[10] ), 
        .B1(n738), .Y(n719) );
  NAND2XL U627 ( .A(curr_time[8]), .B(n724), .Y(n720) );
  AOI211XL U628 ( .A0(n521), .A1(n722), .B0(n530), .C0(n516), .Y(n683) );
  NAND2XL U629 ( .A(n477), .B(curr_time[8]), .Y(n722) );
  NOR2XL U630 ( .A(n666), .B(n678), .Y(n661) );
  NAND2XL U631 ( .A(curr_time[4]), .B(curr_time[3]), .Y(n678) );
  NAND3XL U632 ( .A(n639), .B(n638), .C(n648), .Y(n345) );
  NAND2XL U633 ( .A(n634), .B(n633), .Y(n635) );
  AOI22XL U634 ( .A0(n647), .A1(\intadd_0/SUM[1] ), .B0(\data_path/si_w[17] ), 
        .B1(n548), .Y(n639) );
  NAND3XL U635 ( .A(n613), .B(n612), .C(n648), .Y(n355) );
  NAND2XL U636 ( .A(n608), .B(n607), .Y(n609) );
  AOI22XL U637 ( .A0(n647), .A1(\intadd_1/SUM[1] ), .B0(\data_path/si_w[9] ), 
        .B1(n548), .Y(n613) );
  NAND3XL U638 ( .A(n588), .B(n587), .C(n648), .Y(n365) );
  NAND2XL U639 ( .A(n583), .B(n582), .Y(n584) );
  AOI22XL U640 ( .A0(n647), .A1(\intadd_2/SUM[1] ), .B0(\data_path/si_w[1] ), 
        .B1(n548), .Y(n588) );
  NAND3XL U641 ( .A(n646), .B(n645), .C(n648), .Y(n342) );
  AOI22XL U642 ( .A0(n658), .A1(\intadd_0/SUM[2] ), .B0(n647), .B1(
        \intadd_0/SUM[4] ), .Y(n645) );
  OAI211XL U643 ( .A0(n660), .A1(n642), .B0(n632), .C0(n648), .Y(n346) );
  OAI21XL U644 ( .A0(IM_D[16]), .A1(n741), .B0(n629), .Y(n631) );
  NAND3XL U645 ( .A(n650), .B(n649), .C(n648), .Y(n341) );
  AOI22XL U646 ( .A0(n658), .A1(\intadd_0/SUM[3] ), .B0(n647), .B1(
        \intadd_0/SUM[5] ), .Y(n649) );
  OAI211XL U647 ( .A0(n660), .A1(n591), .B0(n581), .C0(n648), .Y(n366) );
  OAI21XL U648 ( .A0(IM_D[0]), .A1(n741), .B0(n629), .Y(n563) );
  OAI211XL U649 ( .A0(n660), .A1(n616), .B0(n606), .C0(n648), .Y(n356) );
  OAI21XL U650 ( .A0(IM_D[8]), .A1(n741), .B0(n629), .Y(n605) );
  AOI211XL U651 ( .A0(n647), .A1(\intadd_2/SUM[5] ), .B0(n657), .C0(n596), .Y(
        n597) );
  AOI211XL U652 ( .A0(n647), .A1(\intadd_1/SUM[5] ), .B0(n657), .C0(n621), .Y(
        n622) );
  AOI211XL U653 ( .A0(n647), .A1(\intadd_2/SUM[3] ), .B0(n657), .C0(n592), .Y(
        n593) );
  AOI211XL U654 ( .A0(n647), .A1(\intadd_2/SUM[4] ), .B0(n657), .C0(n594), .Y(
        n595) );
  AOI211XL U655 ( .A0(n647), .A1(\intadd_1/SUM[3] ), .B0(n657), .C0(n617), .Y(
        n618) );
  AOI211XL U656 ( .A0(n647), .A1(\intadd_1/SUM[4] ), .B0(n657), .C0(n619), .Y(
        n620) );
  AOI211XL U657 ( .A0(n647), .A1(\intadd_0/SUM[3] ), .B0(n657), .C0(n643), .Y(
        n644) );
  AOI211XL U658 ( .A0(n658), .A1(\intadd_0/SUM[5] ), .B0(n657), .C0(n656), .Y(
        n659) );
  NAND2XL U659 ( .A(\intadd_0/CO ), .B(im_d_w[28]), .Y(n654) );
  AOI211XL U660 ( .A0(n548), .A1(\data_path/si_w[22] ), .B0(n657), .C0(n651), 
        .Y(n652) );
  AOI211XL U661 ( .A0(n647), .A1(\intadd_1/SUM[2] ), .B0(n657), .C0(n614), .Y(
        n615) );
  INVXL U662 ( .A(\intadd_1/SUM[0] ), .Y(n616) );
  AOI211XL U663 ( .A0(\data_path/si_w[6] ), .A1(n548), .B0(n657), .C0(n598), 
        .Y(n599) );
  AOI211XL U664 ( .A0(n647), .A1(\intadd_2/SUM[2] ), .B0(n657), .C0(n589), .Y(
        n590) );
  INVXL U665 ( .A(\intadd_2/SUM[0] ), .Y(n591) );
  AOI211XL U666 ( .A0(n647), .A1(\intadd_0/SUM[2] ), .B0(n657), .C0(n640), .Y(
        n641) );
  INVXL U667 ( .A(\intadd_0/SUM[0] ), .Y(n642) );
  NAND2XL U668 ( .A(n528), .B(n628), .Y(n634) );
  AOI211XL U669 ( .A0(n658), .A1(\intadd_1/SUM[4] ), .B0(n657), .C0(n623), .Y(
        n624) );
  AOI211XL U670 ( .A0(n658), .A1(\intadd_2/SUM[5] ), .B0(n657), .C0(n602), .Y(
        n603) );
  NAND2XL U671 ( .A(\intadd_2/CO ), .B(im_d_w_8), .Y(n601) );
  NAND2XL U672 ( .A(n745), .B(n553), .Y(n583) );
  AOI211XL U673 ( .A0(n658), .A1(\intadd_1/SUM[5] ), .B0(n657), .C0(n626), .Y(
        n627) );
  NOR3XL U674 ( .A(n740), .B(so_mux_sel[0]), .C(so_mux_sel[1]), .Y(n655) );
  AOI211XL U675 ( .A0(expand_sel[3]), .A1(n576), .B0(so_mux_sel[0]), .C0(n575), 
        .Y(n579) );
  NAND2XL U676 ( .A(so_mux_sel[1]), .B(en_so), .Y(n575) );
  AOI31XL U677 ( .A0(expand_sel[2]), .A1(n569), .A2(n568), .B0(n567), .Y(n580)
         );
  AOI211XL U678 ( .A0(n577), .A1(\data_path/si_w[12] ), .B0(expand_sel[2]), 
        .C0(n566), .Y(n567) );
  NAND2XL U679 ( .A(expand_sel[0]), .B(n573), .Y(n565) );
  INVXL U680 ( .A(n769), .Y(n768) );
  AOI222XL U681 ( .A0(n744), .A1(\data_path/si_w[2] ), .B0(n549), .B1(IM_Q[2]), 
        .C0(n731), .C1(CR_Q[2]), .Y(n314) );
  AOI222XL U682 ( .A0(n550), .A1(\data_path/si_w[4] ), .B0(n549), .B1(IM_Q[4]), 
        .C0(n731), .C1(CR_Q[4]), .Y(n313) );
  AOI222XL U683 ( .A0(n550), .A1(\data_path/si_w[8] ), .B0(n549), .B1(IM_Q[8]), 
        .C0(n731), .C1(CR_Q[8]), .Y(n312) );
  AOI222XL U684 ( .A0(n550), .A1(\data_path/si_w[1] ), .B0(n731), .B1(CR_Q[1]), 
        .C0(IM_Q[1]), .C1(n549), .Y(n315) );
  AOI222XL U685 ( .A0(n550), .A1(\data_path/si_w[12] ), .B0(n549), .B1(
        IM_Q[12]), .C0(n731), .C1(CR_Q[12]), .Y(n732) );
  AOI222XL U686 ( .A0(n550), .A1(\data_path/si_w[0] ), .B0(n549), .B1(IM_Q[0]), 
        .C0(n731), .C1(CR_Q[0]), .Y(n555) );
  AOI222XL U687 ( .A0(n550), .A1(\data_path/si_w[10] ), .B0(n549), .B1(
        IM_Q[10]), .C0(n731), .C1(CR_Q[10]), .Y(n721) );
  AOI222XL U688 ( .A0(n550), .A1(\data_path/si_w[11] ), .B0(n549), .B1(
        IM_Q[11]), .C0(n731), .C1(CR_Q[11]), .Y(n726) );
  AOI222XL U689 ( .A0(n550), .A1(\data_path/si_w[7] ), .B0(n549), .B1(IM_Q[7]), 
        .C0(n731), .C1(CR_Q[7]), .Y(n712) );
  AOI222XL U690 ( .A0(n550), .A1(\data_path/si_w[5] ), .B0(n549), .B1(IM_Q[5]), 
        .C0(n731), .C1(CR_Q[5]), .Y(n710) );
  AOI222XL U691 ( .A0(n550), .A1(\data_path/si_w[6] ), .B0(n549), .B1(IM_Q[6]), 
        .C0(n731), .C1(CR_Q[6]), .Y(n711) );
  AOI222XL U692 ( .A0(n550), .A1(\data_path/si_w[3] ), .B0(n549), .B1(IM_Q[3]), 
        .C0(n731), .C1(CR_Q[3]), .Y(n709) );
  AOI222XL U693 ( .A0(n550), .A1(\data_path/si_w[9] ), .B0(n549), .B1(IM_Q[9]), 
        .C0(n731), .C1(CR_Q[9]), .Y(n716) );
  AND2X2 U694 ( .A(si_sel), .B(en_si), .Y(n731) );
  OAI22XL U695 ( .A0(en_photo_num), .A1(n10), .B0(n747), .B1(n746), .Y(n21) );
  NOR3XL U696 ( .A(\data_path/si_w[9] ), .B(\data_path/si_w[0] ), .C(
        \data_path/si_w[3] ), .Y(n557) );
  OA22X1 U697 ( .A0(n551), .A1(\data_path/si_w[2] ), .B0(n473), .B1(
        curr_photo_addr[2]), .Y(n17) );
  OA22X1 U698 ( .A0(n551), .A1(\data_path/si_w[4] ), .B0(n473), .B1(
        curr_photo_addr[4]), .Y(n15) );
  OA22X1 U699 ( .A0(n552), .A1(\data_path/si_w[2] ), .B0(n474), .B1(fb_addr[2]), .Y(n18) );
  OA22X1 U700 ( .A0(n552), .A1(\data_path/si_w[4] ), .B0(n474), .B1(fb_addr[4]), .Y(n16) );
  NAND4XL U701 ( .A(n514), .B(n517), .C(n524), .D(n534), .Y(n556) );
  NOR3XL U702 ( .A(\data_path/si_w[0] ), .B(\data_path/si_w[3] ), .C(n527), 
        .Y(n560) );
  AOI222XL U703 ( .A0(n684), .A1(curr_time[2]), .B0(n738), .B1(
        \data_path/si_w[2] ), .C0(n667), .C1(n669), .Y(n144) );
  AOI222XL U704 ( .A0(\data_path/si_w[5] ), .A1(n738), .B0(curr_time[5]), .B1(
        n737), .C0(n680), .C1(n679), .Y(n681) );
  OAI222XL U705 ( .A0(n523), .A1(n736), .B0(n545), .B1(n735), .C0(n734), .C1(
        n733), .Y(n326) );
  OAI21XL U706 ( .A0(n727), .A1(n516), .B0(n725), .Y(n328) );
  AOI222XL U707 ( .A0(n704), .A1(curr_time[20]), .B0(curr_time[19]), .B1(n703), 
        .C0(n738), .C1(\data_path/si_w[20] ), .Y(n705) );
  OAI31XL U708 ( .A0(curr_time[12]), .A1(n516), .A2(n733), .B0(n730), .Y(n327)
         );
  OAI31XL U709 ( .A0(curr_time[10]), .A1(n539), .A2(n720), .B0(n719), .Y(n329)
         );
  OAI2BB2XL U710 ( .B0(n742), .B1(n741), .A0N(im_d_w_19), .A1N(n740), .Y(n347)
         );
  OAI2BB2XL U711 ( .B0(n715), .B1(n741), .A0N(im_d_w_9), .A1N(n740), .Y(n357)
         );
  NAND2X1 U712 ( .A(\data_path/si_w[0] ), .B(IM_D[0]), .Y(n553) );
  NAND2X2 U713 ( .A(en_so), .B(n554), .Y(n741) );
  OAI2BB1X1 U714 ( .A0N(n583), .A1N(IM_D[1]), .B0(n582), .Y(\intadd_2/CI ) );
  AO22X1 U715 ( .A0(\data_path/si_w[16] ), .A1(n744), .B0(n549), .B1(IM_Q[16]), 
        .Y(n418) );
  AOI2BB2X1 U716 ( .B0(n474), .B1(n531), .A0N(n474), .A1N(fb_addr[0]), .Y(n416) );
  AOI2BB2X1 U717 ( .B0(n473), .B1(n531), .A0N(n473), .A1N(curr_photo_addr[0]), 
        .Y(n415) );
  AOI2BB2X1 U718 ( .B0(n474), .B1(n537), .A0N(n474), .A1N(fb_addr[3]), .Y(n413) );
  AOI2BB2X1 U719 ( .B0(n473), .B1(n537), .A0N(n473), .A1N(curr_photo_addr[3]), 
        .Y(n412) );
  AOI2BB2X1 U720 ( .B0(n474), .B1(n524), .A0N(n474), .A1N(fb_addr[5]), .Y(n410) );
  AOI2BB2X1 U721 ( .B0(n473), .B1(n524), .A0N(n473), .A1N(curr_photo_addr[5]), 
        .Y(n409) );
  AOI2BB2X1 U722 ( .B0(n474), .B1(n534), .A0N(n474), .A1N(fb_addr[6]), .Y(n407) );
  AOI2BB2X1 U723 ( .B0(n473), .B1(n534), .A0N(n473), .A1N(curr_photo_addr[6]), 
        .Y(n406) );
  AOI2BB2X1 U724 ( .B0(n474), .B1(n536), .A0N(n474), .A1N(fb_addr[7]), .Y(n404) );
  AOI2BB2X1 U725 ( .B0(n473), .B1(n536), .A0N(n473), .A1N(curr_photo_addr[7]), 
        .Y(n403) );
  AOI2BB2X1 U726 ( .B0(en_photo_num), .B1(\data_path/si_w[0] ), .A0N(
        en_photo_num), .A1N(photo_num[0]), .Y(n367) );
  OAI21XL U727 ( .A0(\data_path/si_w[0] ), .A1(n707), .B0(en_so), .Y(n562) );
  AOI22X1 U728 ( .A0(\data_path/si_w[0] ), .A1(n563), .B0(IM_D[0]), .B1(n562), 
        .Y(n581) );
  OAI221XL U729 ( .A0(expand_sel[0]), .A1(\data_path/si_w[6] ), .B0(n570), 
        .B1(\data_path/si_w[5] ), .C0(expand_sel[1]), .Y(n568) );
  OAI22XL U730 ( .A0(expand_sel[0]), .A1(\data_path/si_w[10] ), .B0(n570), 
        .B1(\data_path/si_w[9] ), .Y(n564) );
  OAI22XL U731 ( .A0(n517), .A1(n565), .B0(n573), .B1(n564), .Y(n566) );
  OAI22XL U732 ( .A0(expand_sel[0]), .A1(\data_path/si_w[2] ), .B0(n570), .B1(
        \data_path/si_w[1] ), .Y(n572) );
  OAI221XL U733 ( .A0(expand_sel[0]), .A1(\data_path/si_w[4] ), .B0(n570), 
        .B1(\data_path/si_w[3] ), .C0(n573), .Y(n571) );
  OAI21XL U734 ( .A0(n573), .A1(n572), .B0(n571), .Y(n574) );
  OAI2BB2XL U735 ( .B0(expand_sel[2]), .B1(n574), .A0N(expand_sel[2]), .A1N(
        n531), .Y(n576) );
  NAND3BX1 U736 ( .AN(n577), .B(expand_sel[3]), .C(expand_sel[2]), .Y(n578) );
  AOI2BB1X1 U737 ( .A0N(n484), .A1N(n584), .B0(n707), .Y(n586) );
  OAI21XL U738 ( .A0(n584), .A1(n740), .B0(n484), .Y(n585) );
  OAI21XL U739 ( .A0(n586), .A1(n740), .B0(n585), .Y(n587) );
  AO22X1 U740 ( .A0(n740), .A1(IM_D[2]), .B0(\data_path/si_w[2] ), .B1(n548), 
        .Y(n589) );
  OAI21XL U741 ( .A0(n741), .A1(n591), .B0(n590), .Y(n364) );
  AO22X1 U742 ( .A0(\data_path/si_w[3] ), .A1(n548), .B0(n740), .B1(IM_D[3]), 
        .Y(n592) );
  OAI2BB1X1 U743 ( .A0N(n658), .A1N(\intadd_2/SUM[1] ), .B0(n593), .Y(n363) );
  AO22X1 U744 ( .A0(\data_path/si_w[4] ), .A1(n548), .B0(n740), .B1(IM_D[4]), 
        .Y(n594) );
  OAI2BB1X1 U745 ( .A0N(n658), .A1N(\intadd_2/SUM[2] ), .B0(n595), .Y(n362) );
  AO22X1 U746 ( .A0(\data_path/si_w[5] ), .A1(n548), .B0(n740), .B1(IM_D[5]), 
        .Y(n596) );
  OAI2BB1X1 U747 ( .A0N(n658), .A1N(\intadd_2/SUM[3] ), .B0(n597), .Y(n361) );
  OAI2BB2XL U748 ( .B0(\intadd_2/CO ), .B1(im_d_w_8), .A0N(\intadd_2/CO ), 
        .A1N(im_d_w_8), .Y(n600) );
  AO22X1 U749 ( .A0(\intadd_2/SUM[4] ), .A1(n658), .B0(IM_D[6]), .B1(n740), 
        .Y(n598) );
  OAI21XL U750 ( .A0(n600), .A1(n660), .B0(n599), .Y(n360) );
  AOI2BB2X1 U751 ( .B0(im_d_w_9), .B1(n601), .A0N(im_d_w_9), .A1N(n601), .Y(
        n715) );
  AO22X1 U752 ( .A0(\data_path/si_w[7] ), .A1(n548), .B0(n740), .B1(IM_D[7]), 
        .Y(n602) );
  OAI21XL U753 ( .A0(n660), .A1(n715), .B0(n603), .Y(n359) );
  OAI2BB1X1 U754 ( .A0N(n608), .A1N(IM_D[9]), .B0(n607), .Y(\intadd_1/CI ) );
  OAI21XL U755 ( .A0(\data_path/si_w[8] ), .A1(n707), .B0(en_so), .Y(n604) );
  AOI2BB1X1 U756 ( .A0N(n480), .A1N(n609), .B0(n707), .Y(n611) );
  OAI21XL U757 ( .A0(n609), .A1(n740), .B0(n480), .Y(n610) );
  OAI21XL U758 ( .A0(n611), .A1(n740), .B0(n610), .Y(n612) );
  AO22X1 U759 ( .A0(\data_path/si_w[10] ), .A1(n548), .B0(n740), .B1(IM_D[10]), 
        .Y(n614) );
  OAI21XL U760 ( .A0(n741), .A1(n616), .B0(n615), .Y(n354) );
  AO22X1 U761 ( .A0(\data_path/si_w[11] ), .A1(n548), .B0(n740), .B1(IM_D[11]), 
        .Y(n617) );
  OAI2BB1X1 U762 ( .A0N(n658), .A1N(\intadd_1/SUM[1] ), .B0(n618), .Y(n353) );
  AO22X1 U763 ( .A0(\data_path/si_w[12] ), .A1(n548), .B0(n740), .B1(IM_D[12]), 
        .Y(n619) );
  OAI2BB1X1 U764 ( .A0N(n658), .A1N(\intadd_1/SUM[2] ), .B0(n620), .Y(n352) );
  AO22X1 U765 ( .A0(\data_path/si_w[13] ), .A1(n548), .B0(n740), .B1(IM_D[13]), 
        .Y(n621) );
  OAI2BB1X1 U766 ( .A0N(n658), .A1N(\intadd_1/SUM[3] ), .B0(n622), .Y(n351) );
  AO22X1 U767 ( .A0(\data_path/si_w[14] ), .A1(n548), .B0(n740), .B1(IM_D[14]), 
        .Y(n623) );
  OAI21XL U768 ( .A0(n660), .A1(n739), .B0(n624), .Y(n350) );
  AOI2BB2X1 U769 ( .B0(im_d_w_19), .B1(n625), .A0N(im_d_w_19), .A1N(n625), .Y(
        n742) );
  AO22X1 U770 ( .A0(\data_path/si_w[15] ), .A1(n548), .B0(n740), .B1(IM_D[15]), 
        .Y(n626) );
  OAI21XL U771 ( .A0(n660), .A1(n742), .B0(n627), .Y(n349) );
  OAI2BB1X1 U772 ( .A0N(n634), .A1N(IM_D[17]), .B0(n633), .Y(\intadd_0/CI ) );
  OAI21XL U773 ( .A0(\data_path/si_w[16] ), .A1(n707), .B0(en_so), .Y(n630) );
  AOI2BB1X1 U774 ( .A0N(n482), .A1N(n635), .B0(n707), .Y(n637) );
  OAI21XL U775 ( .A0(n635), .A1(n740), .B0(n482), .Y(n636) );
  OAI21XL U776 ( .A0(n637), .A1(n740), .B0(n636), .Y(n638) );
  AO22X1 U777 ( .A0(\data_path/si_w[18] ), .A1(n548), .B0(n740), .B1(IM_D[18]), 
        .Y(n640) );
  OAI21XL U778 ( .A0(n741), .A1(n642), .B0(n641), .Y(n344) );
  AO22X1 U779 ( .A0(\data_path/si_w[19] ), .A1(n548), .B0(n740), .B1(n793), 
        .Y(n643) );
  OAI2BB1X1 U780 ( .A0N(n658), .A1N(\intadd_0/SUM[1] ), .B0(n644), .Y(n343) );
  OAI2BB2XL U781 ( .B0(\intadd_0/CO ), .B1(im_d_w[28]), .A0N(\intadd_0/CO ), 
        .A1N(im_d_w[28]), .Y(n653) );
  AO22X1 U782 ( .A0(\intadd_0/SUM[4] ), .A1(n658), .B0(n790), .B1(n740), .Y(
        n651) );
  OAI21XL U783 ( .A0(n653), .A1(n660), .B0(n652), .Y(n340) );
  AOI2BB2X1 U784 ( .B0(im_d_w[29]), .B1(n654), .A0N(im_d_w[29]), .A1N(n654), 
        .Y(n708) );
  AO22X1 U785 ( .A0(\data_path/si_w[23] ), .A1(n548), .B0(n789), .B1(n740), 
        .Y(n656) );
  OAI21XL U786 ( .A0(n660), .A1(n708), .B0(n659), .Y(n339) );
  OAI22XL U787 ( .A0(curr_time[0]), .A1(n663), .B0(n529), .B1(n684), .Y(n662)
         );
  OAI21XL U788 ( .A0(n736), .A1(n531), .B0(n662), .Y(n336) );
  OAI22XL U789 ( .A0(en_init_time), .A1(n515), .B0(n736), .B1(n745), .Y(n664)
         );
  OAI21XL U790 ( .A0(n736), .A1(n537), .B0(n670), .Y(n335) );
  AO22X1 U791 ( .A0(n738), .A1(\data_path/si_w[6] ), .B0(n684), .B1(
        curr_time[6]), .Y(n333) );
  AO22X1 U792 ( .A0(n738), .A1(\data_path/si_w[7] ), .B0(n684), .B1(
        curr_time[7]), .Y(n332) );
  OAI21XL U793 ( .A0(n736), .A1(n520), .B0(n685), .Y(n331) );
  AOI2BB2X1 U794 ( .B0(n738), .B1(\data_path/si_w[16] ), .A0N(curr_time[16]), 
        .A1N(n699), .Y(n691) );
  OAI21XL U795 ( .A0(n735), .A1(n518), .B0(n691), .Y(n323) );
  OAI22XL U796 ( .A0(curr_time[17]), .A1(n694), .B0(n532), .B1(n695), .Y(n693)
         );
  OAI21XL U797 ( .A0(n736), .A1(n528), .B0(n693), .Y(n322) );
  OAI21XL U798 ( .A0(n696), .A1(n695), .B0(curr_time[18]), .Y(n697) );
  OAI22XL U799 ( .A0(curr_time[19]), .A1(n703), .B0(n546), .B1(n704), .Y(n702)
         );
  OAI21XL U800 ( .A0(n736), .A1(n538), .B0(n702), .Y(n320) );
  AO22X1 U801 ( .A0(n738), .A1(\data_path/si_w[21] ), .B0(n706), .B1(
        curr_time[21]), .Y(n318) );
  AO22X1 U802 ( .A0(n706), .A1(curr_time[22]), .B0(n738), .B1(
        \data_path/si_w[22] ), .Y(n317) );
  OAI22XL U803 ( .A0(n735), .A1(n519), .B0(n736), .B1(n526), .Y(n316) );
  OAI2BB2XL U804 ( .B0(n708), .B1(n741), .A0N(im_d_w[29]), .A1N(n740), .Y(n337) );
  AOI2BB2X1 U805 ( .B0(\data_path/si_w[9] ), .B1(n738), .A0N(n477), .A1N(n720), 
        .Y(n714) );
  OAI21XL U806 ( .A0(n717), .A1(n539), .B0(n714), .Y(n330) );
  AOI2BB2X1 U807 ( .B0(n473), .B1(n527), .A0N(n473), .A1N(curr_photo_addr[9]), 
        .Y(n400) );
  AOI2BB2X1 U808 ( .B0(n474), .B1(n527), .A0N(n474), .A1N(fb_addr[9]), .Y(n401) );
  OAI21XL U809 ( .A0(n477), .A1(n728), .B0(n717), .Y(n718) );
  AOI2BB2X1 U810 ( .B0(n473), .B1(n514), .A0N(n473), .A1N(curr_photo_addr[10]), 
        .Y(n397) );
  AOI2BB2X1 U811 ( .B0(n474), .B1(n514), .A0N(n474), .A1N(fb_addr[10]), .Y(
        n398) );
  AOI2BB1X1 U812 ( .A0N(n723), .A1N(n728), .B0(n737), .Y(n727) );
  AOI2BB2X1 U813 ( .B0(\data_path/si_w[11] ), .B1(n738), .A0N(curr_time[11]), 
        .A1N(n733), .Y(n725) );
  AOI2BB2X1 U814 ( .B0(n473), .B1(n517), .A0N(n473), .A1N(curr_photo_addr[11]), 
        .Y(n394) );
  AOI2BB2X1 U815 ( .B0(n474), .B1(n517), .A0N(n474), .A1N(fb_addr[11]), .Y(
        n395) );
  OAI21XL U816 ( .A0(curr_time[11]), .A1(n728), .B0(n727), .Y(n729) );
  AOI2BB2X1 U817 ( .B0(n473), .B1(n533), .A0N(n473), .A1N(curr_photo_addr[12]), 
        .Y(n391) );
  AOI2BB2X1 U818 ( .B0(n474), .B1(n533), .A0N(n474), .A1N(fb_addr[12]), .Y(
        n392) );
  AOI2BB2X1 U819 ( .B0(n473), .B1(n523), .A0N(n473), .A1N(curr_photo_addr[13]), 
        .Y(n388) );
  AOI2BB2X1 U820 ( .B0(n474), .B1(n523), .A0N(n474), .A1N(fb_addr[13]), .Y(
        n389) );
  AO22X1 U821 ( .A0(\data_path/si_w[13] ), .A1(n744), .B0(n549), .B1(IM_Q[13]), 
        .Y(n390) );
  AO22X1 U822 ( .A0(n738), .A1(\data_path/si_w[14] ), .B0(n737), .B1(
        curr_time[14]), .Y(n325) );
  AOI2BB2X1 U823 ( .B0(n473), .B1(n541), .A0N(n473), .A1N(curr_photo_addr[14]), 
        .Y(n385) );
  AOI2BB2X1 U824 ( .B0(n474), .B1(n541), .A0N(n474), .A1N(fb_addr[14]), .Y(
        n386) );
  AO22X1 U825 ( .A0(\data_path/si_w[14] ), .A1(n744), .B0(n549), .B1(IM_Q[14]), 
        .Y(n387) );
  AO22X1 U826 ( .A0(n738), .A1(\data_path/si_w[15] ), .B0(n737), .B1(
        curr_time[15]), .Y(n324) );
  AOI2BB2X1 U827 ( .B0(n473), .B1(n542), .A0N(n473), .A1N(curr_photo_addr[15]), 
        .Y(n382) );
  AOI2BB2X1 U828 ( .B0(n474), .B1(n542), .A0N(n474), .A1N(fb_addr[15]), .Y(
        n383) );
  AO22X1 U829 ( .A0(\data_path/si_w[15] ), .A1(n744), .B0(n549), .B1(IM_Q[15]), 
        .Y(n384) );
  AOI2BB2X1 U830 ( .B0(n473), .B1(n528), .A0N(n473), .A1N(curr_photo_addr[17]), 
        .Y(n379) );
  AOI2BB2X1 U831 ( .B0(n474), .B1(n528), .A0N(n474), .A1N(fb_addr[17]), .Y(
        n380) );
  AO22X1 U832 ( .A0(\data_path/si_w[17] ), .A1(n744), .B0(n549), .B1(IM_Q[17]), 
        .Y(n381) );
  OAI2BB2XL U833 ( .B0(n739), .B1(n741), .A0N(n740), .A1N(im_d_w_18), .Y(n348)
         );
  AOI2BB2X1 U834 ( .B0(n473), .B1(n535), .A0N(n473), .A1N(curr_photo_addr[18]), 
        .Y(n376) );
  AOI2BB2X1 U835 ( .B0(n474), .B1(n535), .A0N(n474), .A1N(fb_addr[18]), .Y(
        n377) );
  AO22X1 U836 ( .A0(\data_path/si_w[18] ), .A1(n744), .B0(n549), .B1(IM_Q[18]), 
        .Y(n378) );
  AOI2BB2X1 U837 ( .B0(n473), .B1(n538), .A0N(n473), .A1N(curr_photo_addr[19]), 
        .Y(n373) );
  AOI2BB2X1 U838 ( .B0(n474), .B1(n538), .A0N(n474), .A1N(fb_addr[19]), .Y(
        n374) );
  AO22X1 U839 ( .A0(\data_path/si_w[19] ), .A1(n744), .B0(n549), .B1(IM_Q[19]), 
        .Y(n375) );
  AO22X1 U840 ( .A0(\data_path/si_w[20] ), .A1(n744), .B0(n549), .B1(IM_Q[20]), 
        .Y(n372) );
  AO22X1 U841 ( .A0(\data_path/si_w[21] ), .A1(n744), .B0(n549), .B1(IM_Q[21]), 
        .Y(n371) );
  AO22X1 U842 ( .A0(\data_path/si_w[22] ), .A1(n744), .B0(n549), .B1(IM_Q[22]), 
        .Y(n370) );
  AO22X1 U843 ( .A0(\data_path/si_w[23] ), .A1(n744), .B0(n549), .B1(IM_Q[23]), 
        .Y(n369) );
  AO22X1 U844 ( .A0(n473), .A1(\data_path/si_w[16] ), .B0(n551), .B1(
        curr_photo_addr[16]), .Y(n11) );
  AO22X1 U845 ( .A0(n474), .A1(\data_path/si_w[16] ), .B0(n552), .B1(
        fb_addr[16]), .Y(n12) );
  AOI2BB2X1 U846 ( .B0(n473), .B1(n520), .A0N(n473), .A1N(curr_photo_addr[8]), 
        .Y(n13) );
  AOI2BB2X1 U847 ( .B0(n474), .B1(n520), .A0N(n474), .A1N(fb_addr[8]), .Y(n14)
         );
  AOI2BB2X1 U848 ( .B0(n473), .B1(n745), .A0N(n473), .A1N(curr_photo_addr[1]), 
        .Y(n19) );
  AOI2BB2X1 U849 ( .B0(n474), .B1(n745), .A0N(n474), .A1N(fb_addr[1]), .Y(n20)
         );
  OAI22XL U850 ( .A0(\data_path/si_w[0] ), .A1(n745), .B0(n531), .B1(
        \data_path/si_w[1] ), .Y(n746) );
  OAI21XL U851 ( .A0(en_curr_photo_size), .A1(n547), .B0(n748), .Y(n23) );
endmodule

