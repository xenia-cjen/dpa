
module CONT ( clk, reset, im_wen_n, cr_a, curr_time, fb_addr, photo_num, 
        curr_photo_addr, curr_photo_size, en_si, en_init_time, en_fb_addr, 
        en_photo_num, en_curr_photo_addr, en_curr_photo_size, en_so, si_sel, 
        init_time_mux_sel, so_mux_sel, expand_sel, \im_a[19]_BAR , 
        \im_a[18]_BAR , \im_a[17]_BAR , \im_a[16]_BAR , \im_a[15]_BAR , 
        \im_a[14]_BAR , \im_a[13]_BAR , \im_a[12]_BAR , \im_a[11]_BAR , 
        \im_a[10]_BAR , \im_a[9]_BAR , \im_a[8]_BAR , \im_a[7]_BAR , 
        \im_a[6]_BAR , \im_a[5]_BAR , \im_a[4]_BAR , \im_a[3]_BAR , 
        \im_a[2]_BAR , \im_a[1]_BAR , \im_a[0]_BAR , \sftr_n[1] , 
        \sftr_n[0]_BAR  );
  output [8:0] cr_a;
  input [23:0] curr_time;
  input [19:0] fb_addr;
  input [1:0] photo_num;
  input [19:0] curr_photo_addr;
  input [1:0] curr_photo_size;
  output [1:0] so_mux_sel;
  output [3:0] expand_sel;
  input clk, reset;
  output im_wen_n, en_si, en_init_time, en_fb_addr, en_photo_num,
         en_curr_photo_addr, en_curr_photo_size, en_so, si_sel,
         init_time_mux_sel, \im_a[19]_BAR , \im_a[18]_BAR , \im_a[17]_BAR ,
         \im_a[16]_BAR , \im_a[15]_BAR , \im_a[14]_BAR , \im_a[13]_BAR ,
         \im_a[12]_BAR , \im_a[11]_BAR , \im_a[10]_BAR , \im_a[9]_BAR ,
         \im_a[8]_BAR , \im_a[7]_BAR , \im_a[6]_BAR , \im_a[5]_BAR ,
         \im_a[4]_BAR , \im_a[3]_BAR , \im_a[2]_BAR , \im_a[1]_BAR ,
         \im_a[0]_BAR , \sftr_n[1] , \sftr_n[0]_BAR ;
  wire   n2878, n2879, n2880, n2881, n2882, n2883, \state[2] ,
         \next_glb_cntr[1] , \next_write_addr_w[0] , \next_cr_y[0] , \h_0[0] ,
         \m_0[0] , \s_1[3] , \s_0[0] , N88, N89, N1138, N1139, N1140, N1141,
         N1142, N1143, N1144, N1145, N1347, N1348, N1349, N1350, N1351, N1352,
         N1353, N1354, N1355, N1356, N1357, N1358, N1359, N1360, N1361, N1362,
         N1363, N1364, N1365, N1366, N1825, N1826, N1827, N196, next_en_si,
         N2250, N2272, N2292, N2294, \C159/DATA3_0 , \C159/DATA3_1 ,
         \C159/DATA3_2 , \C159/DATA3_3 , \C159/DATA3_4 , \C159/DATA3_5 ,
         \C159/DATA3_6 , \C159/DATA3_7 , \C159/DATA3_8 , \C159/DATA3_9 ,
         \C159/DATA3_10 , \C159/DATA3_11 , \C159/DATA3_12 , \C159/DATA3_13 ,
         \C159/DATA3_14 , \C159/DATA3_15 , \C159/DATA3_16 , \C159/DATA3_17 ,
         \C159/DATA3_18 , \C159/DATA3_19 , \C158/DATA2_7 , \C158/DATA2_8 ,
         \C158/DATA2_9 , \C158/DATA2_10 , \C158/DATA2_11 , \C158/DATA2_12 ,
         \C158/DATA2_13 , \C158/DATA2_14 , \C158/DATA2_15 , \C158/DATA2_16 ,
         \C158/DATA2_17 , n17, n26, n27, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n472, n473, n475, n476, n477, n478, n479,
         n480, n481, n482, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n497, n498, n499, n500, \DP_OP_589J1_125_1438/n26 ,
         \DP_OP_589J1_125_1438/n25 , \C1/Z_19 , \C1/Z_18 , \C1/Z_17 ,
         \C1/Z_16 , \C1/Z_15 , \C1/Z_14 , \C1/Z_13 , \C1/Z_12 , \C1/Z_11 ,
         \C1/Z_10 , \C1/Z_9 , \C1/Z_8 , \C2/Z_19 , \C2/Z_18 , \C2/Z_17 ,
         \C2/Z_16 , \C2/Z_15 , \C2/Z_14 , \C2/Z_13 , \C2/Z_12 , \C2/Z_11 ,
         \C2/Z_10 , \C2/Z_9 , \C2/Z_8 , \C2/Z_7 , \C2/Z_6 , \C2/Z_5 , \C2/Z_4 ,
         \C2/Z_3 , \C2/Z_2 , \C2/Z_1 , \C1/Z_7 , \C1/Z_3 , \C1/Z_2 , \C1/Z_1 ,
         \C1/Z_0 , \DP_OP_229J1_126_7015/I2 , \DP_OP_229J1_126_7015/I3 ,
         \DP_OP_229J1_126_7015/n27 , \DP_OP_229J1_126_7015/n26 ,
         \DP_OP_229J1_126_7015/n25 , \DP_OP_229J1_126_7015/n24 ,
         \DP_OP_229J1_126_7015/n23 , \DP_OP_229J1_126_7015/n21 ,
         \DP_OP_229J1_126_7015/n17 , \DP_OP_229J1_126_7015/n16 ,
         \DP_OP_229J1_126_7015/n8 , \DP_OP_229J1_126_7015/n7 ,
         \DP_OP_229J1_126_7015/n6 , \DP_OP_229J1_126_7015/n5 ,
         \DP_OP_229J1_126_7015/n4 , \DP_OP_229J1_126_7015/n3 ,
         \DP_OP_229J1_126_7015/n2 , \DP_OP_229J1_126_7015/n1 ,
         \DP_OP_559J1_134_6328/n10 , \DP_OP_559J1_134_6328/n9 ,
         \DP_OP_559J1_134_6328/n8 , \DP_OP_559J1_134_6328/n7 ,
         \DP_OP_559J1_134_6328/n6 , \DP_OP_559J1_134_6328/n5 ,
         \DP_OP_559J1_134_6328/n4 , \DP_OP_559J1_134_6328/n3 ,
         \DP_OP_559J1_134_6328/n2 , \DP_OP_559J1_134_6328/n1 ,
         \DP_OP_590J1_137_6981/I5 , \DP_OP_590J1_137_6981/n64 ,
         \DP_OP_590J1_137_6981/n63 , \DP_OP_590J1_137_6981/n62 ,
         \DP_OP_590J1_137_6981/n61 , \DP_OP_590J1_137_6981/n60 ,
         \DP_OP_590J1_137_6981/n59 , \DP_OP_590J1_137_6981/n58 ,
         \DP_OP_590J1_137_6981/n57 , \DP_OP_590J1_137_6981/n56 ,
         \DP_OP_590J1_137_6981/n55 , \DP_OP_590J1_137_6981/n54 ,
         \DP_OP_590J1_137_6981/n53 , \DP_OP_590J1_137_6981/n52 ,
         \DP_OP_590J1_137_6981/n51 , \DP_OP_590J1_137_6981/n50 ,
         \DP_OP_590J1_137_6981/n49 , \DP_OP_590J1_137_6981/n48 ,
         \DP_OP_590J1_137_6981/n47 , \DP_OP_590J1_137_6981/n46 ,
         \DP_OP_590J1_137_6981/n40 , \DP_OP_590J1_137_6981/n39 ,
         \DP_OP_590J1_137_6981/n38 , \DP_OP_590J1_137_6981/n37 ,
         \DP_OP_590J1_137_6981/n36 , \DP_OP_590J1_137_6981/n35 ,
         \DP_OP_590J1_137_6981/n34 , \DP_OP_590J1_137_6981/n33 ,
         \DP_OP_590J1_137_6981/n32 , \DP_OP_590J1_137_6981/n31 ,
         \DP_OP_590J1_137_6981/n30 , \DP_OP_590J1_137_6981/n29 ,
         \DP_OP_590J1_137_6981/n28 , \DP_OP_590J1_137_6981/n27 ,
         \DP_OP_590J1_137_6981/n26 , \DP_OP_590J1_137_6981/n25 ,
         \DP_OP_590J1_137_6981/n24 , \DP_OP_590J1_137_6981/n23 ,
         \DP_OP_590J1_137_6981/n22 , \DP_OP_590J1_137_6981/n20 ,
         \DP_OP_590J1_137_6981/n19 , \DP_OP_590J1_137_6981/n18 ,
         \DP_OP_590J1_137_6981/n17 , \DP_OP_590J1_137_6981/n16 ,
         \DP_OP_590J1_137_6981/n15 , \DP_OP_590J1_137_6981/n14 ,
         \DP_OP_590J1_137_6981/n13 , \DP_OP_590J1_137_6981/n12 ,
         \DP_OP_590J1_137_6981/n11 , \DP_OP_590J1_137_6981/n10 ,
         \DP_OP_590J1_137_6981/n9 , \DP_OP_590J1_137_6981/n8 ,
         \DP_OP_590J1_137_6981/n7 , \DP_OP_590J1_137_6981/n6 ,
         \DP_OP_590J1_137_6981/n5 , \DP_OP_590J1_137_6981/n4 ,
         \DP_OP_590J1_137_6981/n3 , \DP_OP_590J1_137_6981/n2 ,
         \DP_OP_590J1_137_6981/n1 , \intadd_3/A[9] , \intadd_3/A[7] ,
         \intadd_3/A[4] , \intadd_3/A[3] , \intadd_3/A[2] , \intadd_3/A[1] ,
         \intadd_3/A[0] , \intadd_3/B[8] , \intadd_3/B[7] , \intadd_3/B[6] ,
         \intadd_3/B[5] , \intadd_3/B[4] , \intadd_3/B[3] , \intadd_3/B[2] ,
         \intadd_3/B[1] , \intadd_3/B[0] , \intadd_3/CI , \intadd_3/SUM[9] ,
         \intadd_3/SUM[8] , \intadd_3/SUM[7] , \intadd_3/SUM[6] ,
         \intadd_3/SUM[5] , \intadd_3/SUM[4] , \intadd_3/SUM[3] ,
         \intadd_3/SUM[2] , \intadd_3/SUM[1] , \intadd_3/SUM[0] ,
         \intadd_3/n10 , \intadd_3/n9 , \intadd_3/n8 , \intadd_3/n7 ,
         \intadd_3/n6 , \intadd_3/n5 , \intadd_3/n4 , \intadd_3/n3 , n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n12, n14, n16, n19, n21, n23, n25,
         n29, n31, n33, n35, n37, n39, n41, n43, n45, n47, n49, n51, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n177,
         n180, n182, n184, n186, n189, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n474, n483, n484, n496, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877;
  wire   [2:0] next_state;
  wire   [19:0] work_cntr;
  wire   [19:0] next_work_cntr;
  wire   [19:0] global_cntr;
  wire   [19:0] write_addr;
  wire   [19:0] write_cntr;
  wire   [8:0] next_cr_x;
  wire   [3:0] m_1;
  wire   [19:0] read_cntr;
  wire   [8:0] cr_read_cntr;
  wire   [1:0] curr_photo;
  wire   [1:0] next_photo;
  assign \h_0[0]  = curr_time[16];
  assign \m_0[0]  = curr_time[8];
  assign \s_0[0]  = curr_time[0];
  assign en_init_time = N2250;
  assign en_curr_photo_addr = N2272;
  assign en_curr_photo_size = N2292;
  assign init_time_mux_sel = N2294;

  DFFSX1 en_si_reg ( .D(next_en_si), .CK(clk), .SN(n133), .Q(en_si) );
  ADDHXL \DP_OP_229J1_126_7015/U16  ( .A(\C1/Z_0 ), .B(\C1/Z_1 ), .CO(
        \DP_OP_229J1_126_7015/n8 ), .S(\DP_OP_229J1_126_7015/n23 ) );
  ADDFXL \DP_OP_229J1_126_7015/U15  ( .A(\C1/Z_2 ), .B(\C1/Z_1 ), .CI(
        \DP_OP_229J1_126_7015/n8 ), .CO(\DP_OP_229J1_126_7015/n7 ), .S(
        \DP_OP_229J1_126_7015/n24 ) );
  ADDFXL \DP_OP_229J1_126_7015/U14  ( .A(\C1/Z_3 ), .B(\C1/Z_2 ), .CI(
        \DP_OP_229J1_126_7015/n7 ), .CO(\DP_OP_229J1_126_7015/n6 ), .S(
        \DP_OP_229J1_126_7015/n25 ) );
  ADDHXL \DP_OP_229J1_126_7015/U13  ( .A(\C1/Z_3 ), .B(
        \DP_OP_229J1_126_7015/n6 ), .CO(\DP_OP_229J1_126_7015/n27 ), .S(
        \DP_OP_229J1_126_7015/n26 ) );
  AO21X1 \DP_OP_229J1_126_7015/U11  ( .A0(\DP_OP_229J1_126_7015/n23 ), .A1(
        n173), .B0(\DP_OP_229J1_126_7015/I2 ), .Y(\DP_OP_229J1_126_7015/n17 )
         );
  ADDHXL \DP_OP_559J1_134_6328/U11  ( .A(write_addr[10]), .B(n260), .CO(
        \DP_OP_559J1_134_6328/n10 ), .S(\C158/DATA2_8 ) );
  ADDHXL \DP_OP_559J1_134_6328/U10  ( .A(write_addr[11]), .B(
        \DP_OP_559J1_134_6328/n10 ), .CO(\DP_OP_559J1_134_6328/n9 ), .S(
        \C158/DATA2_9 ) );
  ADDHXL \DP_OP_559J1_134_6328/U9  ( .A(write_addr[12]), .B(
        \DP_OP_559J1_134_6328/n9 ), .CO(\DP_OP_559J1_134_6328/n8 ), .S(
        \C158/DATA2_10 ) );
  ADDHXL \DP_OP_559J1_134_6328/U8  ( .A(write_addr[13]), .B(
        \DP_OP_559J1_134_6328/n8 ), .CO(\DP_OP_559J1_134_6328/n7 ), .S(
        \C158/DATA2_11 ) );
  ADDHXL \DP_OP_559J1_134_6328/U7  ( .A(write_addr[14]), .B(
        \DP_OP_559J1_134_6328/n7 ), .CO(\DP_OP_559J1_134_6328/n6 ), .S(
        \C158/DATA2_12 ) );
  ADDHXL \DP_OP_559J1_134_6328/U6  ( .A(write_addr[15]), .B(
        \DP_OP_559J1_134_6328/n6 ), .CO(\DP_OP_559J1_134_6328/n5 ), .S(
        \C158/DATA2_13 ) );
  ADDHXL \DP_OP_559J1_134_6328/U5  ( .A(write_addr[16]), .B(
        \DP_OP_559J1_134_6328/n5 ), .CO(\DP_OP_559J1_134_6328/n4 ), .S(
        \C158/DATA2_14 ) );
  ADDHXL \DP_OP_559J1_134_6328/U4  ( .A(write_addr[17]), .B(
        \DP_OP_559J1_134_6328/n4 ), .CO(\DP_OP_559J1_134_6328/n3 ), .S(
        \C158/DATA2_15 ) );
  ADDHXL \DP_OP_559J1_134_6328/U3  ( .A(write_addr[18]), .B(
        \DP_OP_559J1_134_6328/n3 ), .CO(\DP_OP_559J1_134_6328/n2 ), .S(
        \C158/DATA2_16 ) );
  ADDHXL \DP_OP_559J1_134_6328/U2  ( .A(write_addr[19]), .B(
        \DP_OP_559J1_134_6328/n2 ), .CO(\DP_OP_559J1_134_6328/n1 ), .S(
        \C158/DATA2_17 ) );
  ADDFXL \DP_OP_590J1_137_6981/U61  ( .A(write_addr[1]), .B(fb_addr[1]), .CI(
        \DP_OP_590J1_137_6981/n40 ), .CO(\DP_OP_590J1_137_6981/n39 ), .S(N1348) );
  ADDFXL \DP_OP_590J1_137_6981/U60  ( .A(write_addr[2]), .B(fb_addr[2]), .CI(
        \DP_OP_590J1_137_6981/n39 ), .CO(\DP_OP_590J1_137_6981/n38 ), .S(N1349) );
  ADDFXL \DP_OP_590J1_137_6981/U59  ( .A(write_addr[3]), .B(fb_addr[3]), .CI(
        \DP_OP_590J1_137_6981/n38 ), .CO(\DP_OP_590J1_137_6981/n37 ), .S(N1350) );
  ADDFXL \DP_OP_590J1_137_6981/U58  ( .A(write_addr[4]), .B(fb_addr[4]), .CI(
        \DP_OP_590J1_137_6981/n37 ), .CO(\DP_OP_590J1_137_6981/n36 ), .S(N1351) );
  ADDFXL \DP_OP_590J1_137_6981/U57  ( .A(write_addr[5]), .B(fb_addr[5]), .CI(
        \DP_OP_590J1_137_6981/n36 ), .CO(\DP_OP_590J1_137_6981/n35 ), .S(N1352) );
  ADDFXL \DP_OP_590J1_137_6981/U56  ( .A(write_addr[6]), .B(fb_addr[6]), .CI(
        \DP_OP_590J1_137_6981/n35 ), .CO(\DP_OP_590J1_137_6981/n34 ), .S(N1353) );
  ADDFXL \DP_OP_590J1_137_6981/U55  ( .A(write_addr[7]), .B(fb_addr[7]), .CI(
        \DP_OP_590J1_137_6981/n34 ), .CO(\DP_OP_590J1_137_6981/n33 ), .S(N1354) );
  ADDFXL \DP_OP_590J1_137_6981/U54  ( .A(write_addr[8]), .B(fb_addr[8]), .CI(
        \DP_OP_590J1_137_6981/n33 ), .CO(\DP_OP_590J1_137_6981/n32 ), .S(N1355) );
  ADDFXL \DP_OP_590J1_137_6981/U53  ( .A(write_addr[9]), .B(fb_addr[9]), .CI(
        \DP_OP_590J1_137_6981/n32 ), .CO(\DP_OP_590J1_137_6981/n31 ), .S(N1356) );
  ADDFXL \DP_OP_590J1_137_6981/U52  ( .A(write_addr[10]), .B(fb_addr[10]), 
        .CI(\DP_OP_590J1_137_6981/n31 ), .CO(\DP_OP_590J1_137_6981/n30 ), .S(
        N1357) );
  ADDFXL \DP_OP_590J1_137_6981/U51  ( .A(write_addr[11]), .B(fb_addr[11]), 
        .CI(\DP_OP_590J1_137_6981/n30 ), .CO(\DP_OP_590J1_137_6981/n29 ), .S(
        N1358) );
  ADDFXL \DP_OP_590J1_137_6981/U50  ( .A(write_addr[12]), .B(fb_addr[12]), 
        .CI(\DP_OP_590J1_137_6981/n29 ), .CO(\DP_OP_590J1_137_6981/n28 ), .S(
        N1359) );
  ADDFXL \DP_OP_590J1_137_6981/U49  ( .A(write_addr[13]), .B(fb_addr[13]), 
        .CI(\DP_OP_590J1_137_6981/n28 ), .CO(\DP_OP_590J1_137_6981/n27 ), .S(
        N1360) );
  ADDFXL \DP_OP_590J1_137_6981/U48  ( .A(write_addr[14]), .B(fb_addr[14]), 
        .CI(\DP_OP_590J1_137_6981/n27 ), .CO(\DP_OP_590J1_137_6981/n26 ), .S(
        N1361) );
  ADDFXL \DP_OP_590J1_137_6981/U47  ( .A(write_addr[15]), .B(fb_addr[15]), 
        .CI(\DP_OP_590J1_137_6981/n26 ), .CO(\DP_OP_590J1_137_6981/n25 ), .S(
        N1362) );
  ADDFXL \DP_OP_590J1_137_6981/U46  ( .A(write_addr[16]), .B(fb_addr[16]), 
        .CI(\DP_OP_590J1_137_6981/n25 ), .CO(\DP_OP_590J1_137_6981/n24 ), .S(
        N1363) );
  ADDFXL \DP_OP_590J1_137_6981/U45  ( .A(write_addr[17]), .B(fb_addr[17]), 
        .CI(\DP_OP_590J1_137_6981/n24 ), .CO(\DP_OP_590J1_137_6981/n23 ), .S(
        N1364) );
  ADDFXL \DP_OP_590J1_137_6981/U44  ( .A(write_addr[18]), .B(fb_addr[18]), 
        .CI(\DP_OP_590J1_137_6981/n23 ), .CO(\DP_OP_590J1_137_6981/n22 ), .S(
        N1365) );
  AO22X1 \DP_OP_590J1_137_6981/U40  ( .A0(N1348), .A1(n312), .B0(
        \DP_OP_590J1_137_6981/I5 ), .B1(\C2/Z_1 ), .Y(
        \DP_OP_590J1_137_6981/n46 ) );
  AO22X1 \DP_OP_590J1_137_6981/U39  ( .A0(N1349), .A1(n312), .B0(
        \DP_OP_590J1_137_6981/I5 ), .B1(\C2/Z_2 ), .Y(
        \DP_OP_590J1_137_6981/n47 ) );
  AO22X1 \DP_OP_590J1_137_6981/U38  ( .A0(N1350), .A1(n312), .B0(
        \DP_OP_590J1_137_6981/I5 ), .B1(\C2/Z_3 ), .Y(
        \DP_OP_590J1_137_6981/n48 ) );
  AO22X1 \DP_OP_590J1_137_6981/U37  ( .A0(N1351), .A1(n312), .B0(
        \DP_OP_590J1_137_6981/I5 ), .B1(\C2/Z_4 ), .Y(
        \DP_OP_590J1_137_6981/n49 ) );
  AO22X1 \DP_OP_590J1_137_6981/U36  ( .A0(N1352), .A1(n312), .B0(
        \DP_OP_590J1_137_6981/I5 ), .B1(\C2/Z_5 ), .Y(
        \DP_OP_590J1_137_6981/n50 ) );
  AO22X1 \DP_OP_590J1_137_6981/U35  ( .A0(N1353), .A1(n312), .B0(
        \DP_OP_590J1_137_6981/I5 ), .B1(\C2/Z_6 ), .Y(
        \DP_OP_590J1_137_6981/n51 ) );
  AO22X1 \DP_OP_590J1_137_6981/U34  ( .A0(N1354), .A1(n312), .B0(
        \DP_OP_590J1_137_6981/I5 ), .B1(\C2/Z_7 ), .Y(
        \DP_OP_590J1_137_6981/n52 ) );
  AO22X1 \DP_OP_590J1_137_6981/U33  ( .A0(N1355), .A1(n312), .B0(
        \DP_OP_590J1_137_6981/I5 ), .B1(\C2/Z_8 ), .Y(
        \DP_OP_590J1_137_6981/n53 ) );
  AO22X1 \DP_OP_590J1_137_6981/U32  ( .A0(N1356), .A1(n312), .B0(
        \DP_OP_590J1_137_6981/I5 ), .B1(\C2/Z_9 ), .Y(
        \DP_OP_590J1_137_6981/n54 ) );
  AO22X1 \DP_OP_590J1_137_6981/U31  ( .A0(N1357), .A1(n312), .B0(
        \DP_OP_590J1_137_6981/I5 ), .B1(\C2/Z_10 ), .Y(
        \DP_OP_590J1_137_6981/n55 ) );
  AO22X1 \DP_OP_590J1_137_6981/U30  ( .A0(N1358), .A1(n312), .B0(
        \DP_OP_590J1_137_6981/I5 ), .B1(\C2/Z_11 ), .Y(
        \DP_OP_590J1_137_6981/n56 ) );
  AO22X1 \DP_OP_590J1_137_6981/U29  ( .A0(N1359), .A1(n312), .B0(
        \DP_OP_590J1_137_6981/I5 ), .B1(\C2/Z_12 ), .Y(
        \DP_OP_590J1_137_6981/n57 ) );
  AO22X1 \DP_OP_590J1_137_6981/U28  ( .A0(N1360), .A1(n312), .B0(
        \DP_OP_590J1_137_6981/I5 ), .B1(\C2/Z_13 ), .Y(
        \DP_OP_590J1_137_6981/n58 ) );
  AO22X1 \DP_OP_590J1_137_6981/U27  ( .A0(N1361), .A1(n312), .B0(
        \DP_OP_590J1_137_6981/I5 ), .B1(\C2/Z_14 ), .Y(
        \DP_OP_590J1_137_6981/n59 ) );
  AO22X1 \DP_OP_590J1_137_6981/U26  ( .A0(N1362), .A1(n312), .B0(
        \DP_OP_590J1_137_6981/I5 ), .B1(\C2/Z_15 ), .Y(
        \DP_OP_590J1_137_6981/n60 ) );
  AO22X1 \DP_OP_590J1_137_6981/U25  ( .A0(N1363), .A1(si_sel), .B0(
        \DP_OP_590J1_137_6981/I5 ), .B1(\C2/Z_16 ), .Y(
        \DP_OP_590J1_137_6981/n61 ) );
  AO22X1 \DP_OP_590J1_137_6981/U24  ( .A0(N1364), .A1(si_sel), .B0(
        \DP_OP_590J1_137_6981/I5 ), .B1(\C2/Z_17 ), .Y(
        \DP_OP_590J1_137_6981/n62 ) );
  AO22X1 \DP_OP_590J1_137_6981/U23  ( .A0(N1365), .A1(si_sel), .B0(
        \DP_OP_590J1_137_6981/I5 ), .B1(\C2/Z_18 ), .Y(
        \DP_OP_590J1_137_6981/n63 ) );
  AO22X1 \DP_OP_590J1_137_6981/U22  ( .A0(N1366), .A1(si_sel), .B0(
        \DP_OP_590J1_137_6981/I5 ), .B1(\C2/Z_19 ), .Y(
        \DP_OP_590J1_137_6981/n64 ) );
  ADDFXL \DP_OP_590J1_137_6981/U20  ( .A(\DP_OP_590J1_137_6981/n20 ), .B(n730), 
        .CI(\DP_OP_590J1_137_6981/n46 ), .CO(\DP_OP_590J1_137_6981/n19 ), .S(
        \C159/DATA3_1 ) );
  ADDFXL \DP_OP_590J1_137_6981/U19  ( .A(\DP_OP_590J1_137_6981/n47 ), .B(n731), 
        .CI(\DP_OP_590J1_137_6981/n19 ), .CO(\DP_OP_590J1_137_6981/n18 ), .S(
        \C159/DATA3_2 ) );
  ADDFXL \DP_OP_590J1_137_6981/U18  ( .A(\DP_OP_590J1_137_6981/n48 ), .B(n732), 
        .CI(\DP_OP_590J1_137_6981/n18 ), .CO(\DP_OP_590J1_137_6981/n17 ), .S(
        \C159/DATA3_3 ) );
  ADDFXL \DP_OP_590J1_137_6981/U17  ( .A(\DP_OP_590J1_137_6981/n49 ), .B(n733), 
        .CI(\DP_OP_590J1_137_6981/n17 ), .CO(\DP_OP_590J1_137_6981/n16 ), .S(
        \C159/DATA3_4 ) );
  ADDFXL \DP_OP_590J1_137_6981/U16  ( .A(\DP_OP_590J1_137_6981/n50 ), .B(n734), 
        .CI(\DP_OP_590J1_137_6981/n16 ), .CO(\DP_OP_590J1_137_6981/n15 ), .S(
        \C159/DATA3_5 ) );
  ADDFXL \DP_OP_590J1_137_6981/U15  ( .A(\DP_OP_590J1_137_6981/n51 ), .B(n735), 
        .CI(\DP_OP_590J1_137_6981/n15 ), .CO(\DP_OP_590J1_137_6981/n14 ), .S(
        \C159/DATA3_6 ) );
  ADDFXL \DP_OP_590J1_137_6981/U14  ( .A(\DP_OP_590J1_137_6981/n52 ), .B(n736), 
        .CI(\DP_OP_590J1_137_6981/n14 ), .CO(\DP_OP_590J1_137_6981/n13 ), .S(
        \C159/DATA3_7 ) );
  ADDFXL \DP_OP_590J1_137_6981/U13  ( .A(\DP_OP_590J1_137_6981/n53 ), .B(
        \C1/Z_8 ), .CI(\DP_OP_590J1_137_6981/n13 ), .CO(
        \DP_OP_590J1_137_6981/n12 ), .S(\C159/DATA3_8 ) );
  ADDFXL \DP_OP_590J1_137_6981/U12  ( .A(\DP_OP_590J1_137_6981/n54 ), .B(
        \C1/Z_9 ), .CI(\DP_OP_590J1_137_6981/n12 ), .CO(
        \DP_OP_590J1_137_6981/n11 ), .S(\C159/DATA3_9 ) );
  ADDFXL \DP_OP_590J1_137_6981/U11  ( .A(\DP_OP_590J1_137_6981/n55 ), .B(
        \C1/Z_10 ), .CI(\DP_OP_590J1_137_6981/n11 ), .CO(
        \DP_OP_590J1_137_6981/n10 ), .S(\C159/DATA3_10 ) );
  ADDFXL \DP_OP_590J1_137_6981/U10  ( .A(\DP_OP_590J1_137_6981/n56 ), .B(
        \C1/Z_11 ), .CI(\DP_OP_590J1_137_6981/n10 ), .CO(
        \DP_OP_590J1_137_6981/n9 ), .S(\C159/DATA3_11 ) );
  ADDFXL \DP_OP_590J1_137_6981/U9  ( .A(\DP_OP_590J1_137_6981/n57 ), .B(
        \C1/Z_12 ), .CI(\DP_OP_590J1_137_6981/n9 ), .CO(
        \DP_OP_590J1_137_6981/n8 ), .S(\C159/DATA3_12 ) );
  ADDFXL \DP_OP_590J1_137_6981/U8  ( .A(\DP_OP_590J1_137_6981/n58 ), .B(
        \C1/Z_13 ), .CI(\DP_OP_590J1_137_6981/n8 ), .CO(
        \DP_OP_590J1_137_6981/n7 ), .S(\C159/DATA3_13 ) );
  ADDFXL \DP_OP_590J1_137_6981/U7  ( .A(\DP_OP_590J1_137_6981/n59 ), .B(
        \C1/Z_14 ), .CI(\DP_OP_590J1_137_6981/n7 ), .CO(
        \DP_OP_590J1_137_6981/n6 ), .S(\C159/DATA3_14 ) );
  ADDFXL \DP_OP_590J1_137_6981/U6  ( .A(\DP_OP_590J1_137_6981/n60 ), .B(
        \C1/Z_15 ), .CI(\DP_OP_590J1_137_6981/n6 ), .CO(
        \DP_OP_590J1_137_6981/n5 ), .S(\C159/DATA3_15 ) );
  ADDFXL \DP_OP_590J1_137_6981/U5  ( .A(\DP_OP_590J1_137_6981/n61 ), .B(
        \C1/Z_16 ), .CI(\DP_OP_590J1_137_6981/n5 ), .CO(
        \DP_OP_590J1_137_6981/n4 ), .S(\C159/DATA3_16 ) );
  ADDFXL \DP_OP_590J1_137_6981/U4  ( .A(\DP_OP_590J1_137_6981/n62 ), .B(
        \C1/Z_17 ), .CI(\DP_OP_590J1_137_6981/n4 ), .CO(
        \DP_OP_590J1_137_6981/n3 ), .S(\C159/DATA3_17 ) );
  ADDFXL \DP_OP_590J1_137_6981/U3  ( .A(\DP_OP_590J1_137_6981/n63 ), .B(
        \C1/Z_18 ), .CI(\DP_OP_590J1_137_6981/n3 ), .CO(
        \DP_OP_590J1_137_6981/n2 ), .S(\C159/DATA3_18 ) );
  ADDFXL \intadd_3/U11  ( .A(\intadd_3/A[0] ), .B(\intadd_3/B[0] ), .CI(
        \intadd_3/CI ), .CO(\intadd_3/n10 ), .S(\intadd_3/SUM[0] ) );
  ADDFXL \intadd_3/U10  ( .A(\intadd_3/A[1] ), .B(\intadd_3/B[1] ), .CI(
        \intadd_3/n10 ), .CO(\intadd_3/n9 ), .S(\intadd_3/SUM[1] ) );
  ADDFXL \intadd_3/U9  ( .A(\intadd_3/A[2] ), .B(\intadd_3/B[2] ), .CI(
        \intadd_3/n9 ), .CO(\intadd_3/n8 ), .S(\intadd_3/SUM[2] ) );
  ADDFXL \intadd_3/U8  ( .A(\intadd_3/A[3] ), .B(\intadd_3/B[3] ), .CI(
        \intadd_3/n8 ), .CO(\intadd_3/n7 ), .S(\intadd_3/SUM[3] ) );
  ADDFXL \intadd_3/U7  ( .A(\intadd_3/A[4] ), .B(\intadd_3/B[4] ), .CI(
        \intadd_3/n7 ), .CO(\intadd_3/n6 ), .S(\intadd_3/SUM[4] ) );
  ADDFXL \intadd_3/U6  ( .A(\DP_OP_589J1_125_1438/n26 ), .B(\intadd_3/B[5] ), 
        .CI(\intadd_3/n6 ), .CO(\intadd_3/n5 ), .S(\intadd_3/SUM[5] ) );
  ADDFXL \intadd_3/U4  ( .A(\intadd_3/A[7] ), .B(\intadd_3/B[7] ), .CI(
        \intadd_3/n4 ), .CO(\intadd_3/n3 ), .S(\intadd_3/SUM[7] ) );
  ADDFXL \intadd_3/U5  ( .A(\DP_OP_589J1_125_1438/n25 ), .B(\intadd_3/B[6] ), 
        .CI(\intadd_3/n5 ), .CO(\intadd_3/n4 ), .S(\intadd_3/SUM[6] ) );
  ADDHXL \DP_OP_229J1_126_7015/U6  ( .A(N88), .B(\DP_OP_229J1_126_7015/n16 ), 
        .CO(\DP_OP_229J1_126_7015/n5 ), .S(N1141) );
  XOR2XL \DP_OP_590J1_137_6981/U2  ( .A(\DP_OP_590J1_137_6981/n64 ), .B(
        \C1/Z_19 ), .Y(\DP_OP_590J1_137_6981/n1 ) );
  XOR2XL \DP_OP_590J1_137_6981/U1  ( .A(\DP_OP_590J1_137_6981/n2 ), .B(
        \DP_OP_590J1_137_6981/n1 ), .Y(\C159/DATA3_19 ) );
  AND2XL \DP_OP_229J1_126_7015/U12  ( .A(\C1/Z_0 ), .B(n173), .Y(
        \DP_OP_229J1_126_7015/n16 ) );
  AND2XL \DP_OP_229J1_126_7015/U7  ( .A(\DP_OP_229J1_126_7015/n27 ), .B(n173), 
        .Y(\DP_OP_229J1_126_7015/n21 ) );
  DFFSX2 \state_reg[0]  ( .D(n17), .CK(clk), .SN(n133), .Q(n27), .QN(n258) );
  ADDHX1 \DP_OP_590J1_137_6981/U62  ( .A(fb_addr[0]), .B(
        \next_write_addr_w[0] ), .CO(\DP_OP_590J1_137_6981/n40 ), .S(N1347) );
  DFFRX2 \global_cntr_reg[1]  ( .D(\next_glb_cntr[1] ), .CK(clk), .RN(n770), 
        .Q(global_cntr[1]), .QN(n290) );
  DFFRX2 \work_cntr_reg[10]  ( .D(next_work_cntr[10]), .CK(clk), .RN(n770), 
        .Q(work_cntr[10]), .QN(n228) );
  DFFRX2 \work_cntr_reg[18]  ( .D(next_work_cntr[18]), .CK(clk), .RN(n770), 
        .Q(work_cntr[18]), .QN(n252) );
  DFFRX2 \work_cntr_reg[3]  ( .D(next_work_cntr[3]), .CK(clk), .RN(n770), .Q(
        N1827), .QN(n273) );
  DFFRX2 \work_cntr_reg[16]  ( .D(next_work_cntr[16]), .CK(clk), .RN(n770), 
        .Q(work_cntr[16]), .QN(n257) );
  DFFRX2 \work_cntr_reg[7]  ( .D(next_work_cntr[7]), .CK(clk), .RN(n770), .Q(
        work_cntr[7]), .QN(n268) );
  DFFRX2 \work_cntr_reg[17]  ( .D(next_work_cntr[17]), .CK(clk), .RN(n770), 
        .Q(work_cntr[17]), .QN(n231) );
  DFFRX2 \work_cntr_reg[9]  ( .D(n136), .CK(clk), .RN(n770), .Q(work_cntr[9]), 
        .QN(n261) );
  DFFRX2 \work_cntr_reg[6]  ( .D(next_work_cntr[6]), .CK(clk), .RN(n770), .Q(
        work_cntr[6]), .QN(n264) );
  DFFRX2 \write_addr_reg/q_reg[14]  ( .D(n439), .CK(clk), .RN(n770), .Q(
        write_addr[14]), .QN(n224) );
  DFFRX2 \write_addr_reg/q_reg[17]  ( .D(n436), .CK(clk), .RN(n770), .Q(
        write_addr[17]), .QN(n283) );
  DFFRX2 \write_addr_reg/q_reg[19]  ( .D(n434), .CK(clk), .RN(n770), .Q(
        write_addr[19]), .QN(n282) );
  DFFRX2 \write_addr_reg/q_reg[15]  ( .D(n438), .CK(clk), .RN(n770), .Q(
        write_addr[15]), .QN(n299) );
  DFFRX2 \write_cntr_reg/q_reg[9]  ( .D(n490), .CK(clk), .RN(n770), .Q(
        write_cntr[9]), .QN(n267) );
  DFFRX2 \write_cntr_reg/q_reg[8]  ( .D(n497), .CK(clk), .RN(n770), .Q(
        write_cntr[8]), .QN(n269) );
  DFFRX2 \write_cntr_reg/q_reg[7]  ( .D(n491), .CK(clk), .RN(n770), .Q(
        write_cntr[7]), .QN(n272) );
  DFFRX2 \write_cntr_reg/q_reg[6]  ( .D(n492), .CK(clk), .RN(n770), .Q(
        write_cntr[6]), .QN(n287) );
  DFFRX2 \write_cntr_reg/q_reg[5]  ( .D(n493), .CK(clk), .RN(n770), .Q(
        write_cntr[5]), .QN(n274) );
  DFFRX2 \write_cntr_reg/q_reg[10]  ( .D(n489), .CK(clk), .RN(n770), .Q(
        write_cntr[10]), .QN(n199) );
  DFFRX2 \write_addr_reg/q_reg[16]  ( .D(n437), .CK(clk), .RN(n770), .Q(
        write_addr[16]), .QN(n280) );
  DFFRX2 \write_addr_reg/q_reg[1]  ( .D(n481), .CK(clk), .RN(n770), .Q(
        write_addr[1]), .QN(n288) );
  DFFRX2 \write_addr_reg/q_reg[2]  ( .D(n480), .CK(clk), .RN(n770), .Q(
        write_addr[2]), .QN(n238) );
  DFFRX2 \write_addr_reg/q_reg[5]  ( .D(n477), .CK(clk), .RN(n770), .Q(
        write_addr[5]), .QN(n293) );
  DFFRX2 \write_addr_reg/q_reg[7]  ( .D(n475), .CK(clk), .RN(n770), .Q(
        write_addr[7]), .QN(n295) );
  DFFRX2 \write_addr_reg/q_reg[9]  ( .D(n444), .CK(clk), .RN(n770), .Q(
        write_addr[9]), .QN(n294) );
  DFFRX2 \write_addr_reg/q_reg[12]  ( .D(n441), .CK(clk), .RN(n770), .Q(
        write_addr[12]), .QN(n297) );
  DFFRX2 \write_addr_reg/q_reg[13]  ( .D(n440), .CK(clk), .RN(n770), .Q(
        write_addr[13]), .QN(n296) );
  DFFRX2 \write_addr_reg/q_reg[11]  ( .D(n442), .CK(clk), .RN(n770), .Q(
        write_addr[11]), .QN(n223) );
  DFFRX2 \read_cntr_reg/q_reg[0]  ( .D(n473), .CK(clk), .RN(n770), .Q(
        read_cntr[0]), .QN(n285) );
  DFFRX1 \global_cntr_reg[0]  ( .D(n253), .CK(clk), .RN(n133), .Q(
        global_cntr[0]), .QN(n253) );
  DFFRX1 \global_cntr_reg[2]  ( .D(n768), .CK(clk), .RN(n315), .Q(
        global_cntr[2]), .QN(n254) );
  DFFRX1 \global_cntr_reg[3]  ( .D(n766), .CK(clk), .RN(n133), .Q(
        global_cntr[3]), .QN(n291) );
  DFFRX1 \global_cntr_reg[4]  ( .D(n765), .CK(clk), .RN(n133), .Q(
        global_cntr[4]), .QN(n242) );
  DFFRX1 \global_cntr_reg[6]  ( .D(n756), .CK(clk), .RN(n315), .Q(
        global_cntr[6]), .QN(n244) );
  DFFRX1 \global_cntr_reg[7]  ( .D(n755), .CK(clk), .RN(n315), .Q(
        global_cntr[7]), .QN(n298) );
  DFFRX1 \global_cntr_reg[8]  ( .D(n754), .CK(clk), .RN(n315), .Q(
        global_cntr[8]), .QN(n243) );
  DFFRX1 \global_cntr_reg[9]  ( .D(n753), .CK(clk), .RN(n770), .Q(
        global_cntr[9]), .QN(n240) );
  DFFRX1 \global_cntr_reg[10]  ( .D(n752), .CK(clk), .RN(n770), .Q(
        global_cntr[10]), .QN(n247) );
  DFFRX1 \global_cntr_reg[11]  ( .D(n763), .CK(clk), .RN(n133), .Q(
        global_cntr[11]), .QN(n300) );
  DFFRX1 \global_cntr_reg[12]  ( .D(n762), .CK(clk), .RN(n315), .Q(
        global_cntr[12]), .QN(n249) );
  DFFRX1 \global_cntr_reg[14]  ( .D(n760), .CK(clk), .RN(n315), .Q(
        global_cntr[14]), .QN(n248) );
  DFFRX1 \global_cntr_reg[16]  ( .D(n757), .CK(clk), .RN(n133), .Q(
        global_cntr[16]), .QN(n250) );
  DFFRX1 \global_cntr_reg[17]  ( .D(n751), .CK(clk), .RN(n770), .Q(
        global_cntr[17]), .QN(n256) );
  DFFRX1 \global_cntr_reg[18]  ( .D(n750), .CK(clk), .RN(n315), .Q(
        global_cntr[18]), .QN(n218) );
  DFFRX1 \state_reg[1]  ( .D(next_state[1]), .CK(clk), .RN(n315), .Q(n255), 
        .QN(n26) );
  DFFRX1 \state_reg[2]  ( .D(next_state[2]), .CK(clk), .RN(n315), .Q(
        \state[2] ), .QN(n229) );
  DFFRX1 \curr_photo_reg[1]  ( .D(next_photo[1]), .CK(clk), .RN(n133), .Q(
        curr_photo[1]), .QN(n304) );
  DFFRX1 \curr_photo_reg[0]  ( .D(next_photo[0]), .CK(clk), .RN(n315), .Q(
        curr_photo[0]), .QN(n305) );
  DFFRX1 \write_addr_reg/q_reg[18]  ( .D(n435), .CK(clk), .RN(n315), .Q(
        write_addr[18]), .QN(n281) );
  DFFRX1 \write_cntr_reg/q_reg[13]  ( .D(n486), .CK(clk), .RN(n133), .Q(
        write_cntr[13]), .QN(n279) );
  DFFRX1 \write_cntr_reg/q_reg[11]  ( .D(n488), .CK(clk), .RN(n133), .Q(
        write_cntr[11]), .QN(n278) );
  DFFRX1 \write_cntr_reg/q_reg[4]  ( .D(n498), .CK(clk), .RN(n315), .Q(
        write_cntr[4]), .QN(n275) );
  DFFRX1 \write_cntr_reg/q_reg[3]  ( .D(n494), .CK(clk), .RN(n315), .Q(
        write_cntr[3]), .QN(n276) );
  DFFRX1 \write_cntr_reg/q_reg[1]  ( .D(n500), .CK(clk), .RN(n133), .Q(
        write_cntr[1]), .QN(n262) );
  DFFRX1 \write_cntr_reg/q_reg[0]  ( .D(n495), .CK(clk), .RN(n133), .Q(
        write_cntr[0]), .QN(n220) );
  DFFRX1 \write_cntr_reg/q_reg[14]  ( .D(n485), .CK(clk), .RN(n133), .Q(
        write_cntr[14]), .QN(n234) );
  DFFRX1 \write_addr_reg/q_reg[0]  ( .D(n482), .CK(clk), .RN(n133), .Q(
        \next_write_addr_w[0] ), .QN(n236) );
  DFFRX1 \write_addr_reg/q_reg[3]  ( .D(n479), .CK(clk), .RN(n315), .Q(
        write_addr[3]), .QN(n289) );
  DFFRX1 \write_addr_reg/q_reg[6]  ( .D(n476), .CK(clk), .RN(n315), .Q(
        write_addr[6]), .QN(n222) );
  DFFRX1 \write_addr_reg/q_reg[10]  ( .D(n443), .CK(clk), .RN(n315), .Q(
        write_addr[10]), .QN(n292) );
  DFFRX1 \read_cntr_reg/q_reg[1]  ( .D(n472), .CK(clk), .RN(n133), .Q(
        read_cntr[1]), .QN(n237) );
  DFFRX1 \cr_read_cntr_reg/q_reg[2]  ( .D(n452), .CK(clk), .RN(n133), .Q(N1140), .QN(n303) );
  DFFRX1 \cr_read_cntr_reg/q_reg[4]  ( .D(n450), .CK(clk), .RN(n133), .Q(
        cr_read_cntr[4]), .QN(n302) );
  DFFRX1 \cr_read_cntr_reg/q_reg[6]  ( .D(n448), .CK(clk), .RN(n133), .Q(
        cr_read_cntr[6]), .QN(n301) );
  DFFRX1 \cr_read_cntr_reg/q_reg[8]  ( .D(n446), .CK(clk), .RN(n315), .Q(
        cr_read_cntr[8]), .QN(n225) );
  DFFRX1 \global_cntr_reg[5]  ( .D(n764), .CK(clk), .RN(n315), .Q(
        global_cntr[5]) );
  DFFRX1 \global_cntr_reg[13]  ( .D(n761), .CK(clk), .RN(n315), .Q(
        global_cntr[13]) );
  DFFRX1 \global_cntr_reg[15]  ( .D(n759), .CK(clk), .RN(n315), .Q(
        global_cntr[15]) );
  DFFRX1 \global_cntr_reg[19]  ( .D(n749), .CK(clk), .RN(n770), .Q(
        global_cntr[19]) );
  DFFRX1 \write_cntr_reg/q_reg[2]  ( .D(n499), .CK(clk), .RN(n770), .Q(
        write_cntr[2]) );
  DFFRX1 \cr_read_cntr_reg/q_reg[0]  ( .D(n454), .CK(clk), .RN(n133), .Q(N1138), .QN(n5) );
  DFFRX1 \cr_read_cntr_reg/q_reg[3]  ( .D(n451), .CK(clk), .RN(n133), .Q(
        cr_read_cntr[3]) );
  DFFRX1 \cr_read_cntr_reg/q_reg[5]  ( .D(n449), .CK(clk), .RN(n770), .Q(
        cr_read_cntr[5]) );
  DFFRX1 \cr_read_cntr_reg/q_reg[1]  ( .D(n453), .CK(clk), .RN(n133), .Q(N1139), .QN(n7) );
  DFFRX1 \cr_read_cntr_reg/q_reg[7]  ( .D(n447), .CK(clk), .RN(n770), .Q(
        cr_read_cntr[7]) );
  DFFRX4 \work_cntr_reg[1]  ( .D(next_work_cntr[1]), .CK(clk), .RN(n770), .Q(
        N1825), .QN(n232) );
  DFFRX4 \work_cntr_reg[14]  ( .D(next_work_cntr[14]), .CK(clk), .RN(n770), 
        .Q(work_cntr[14]), .QN(n216) );
  DFFRX4 \work_cntr_reg[4]  ( .D(next_work_cntr[4]), .CK(clk), .RN(n770), .Q(
        work_cntr[4]), .QN(n270) );
  DFFRX4 \work_cntr_reg[13]  ( .D(next_work_cntr[13]), .CK(clk), .RN(n770), 
        .Q(work_cntr[13]), .QN(n2423) );
  DFFRX4 \work_cntr_reg[12]  ( .D(next_work_cntr[12]), .CK(clk), .RN(n770), 
        .Q(work_cntr[12]), .QN(n217) );
  DFFRX4 \work_cntr_reg[2]  ( .D(next_work_cntr[2]), .CK(clk), .RN(n770), .Q(
        N1826), .QN(n263) );
  DFFRX4 \work_cntr_reg[5]  ( .D(n2224), .CK(clk), .RN(n770), .Q(work_cntr[5]), 
        .QN(n221) );
  DFFRX4 \work_cntr_reg[19]  ( .D(next_work_cntr[19]), .CK(clk), .RN(n770), 
        .Q(work_cntr[19]), .QN(n259) );
  DFFRX2 \write_addr_reg/q_reg[4]  ( .D(n478), .CK(clk), .RN(n315), .Q(
        write_addr[4]), .QN(n741) );
  DFFRX4 \work_cntr_reg[0]  ( .D(next_work_cntr[0]), .CK(clk), .RN(n770), .Q(
        N196), .QN(n284) );
  DFFRX4 \work_cntr_reg[15]  ( .D(next_work_cntr[15]), .CK(clk), .RN(n770), 
        .Q(work_cntr[15]), .QN(n227) );
  DFFRX4 \write_addr_reg/q_reg[8]  ( .D(n445), .CK(clk), .RN(n770), .Q(
        write_addr[8]), .QN(n235) );
  DFFRX4 \work_cntr_reg[8]  ( .D(next_work_cntr[8]), .CK(clk), .RN(n770), .Q(
        work_cntr[8]), .QN(n266) );
  DFFRX4 \work_cntr_reg[11]  ( .D(next_work_cntr[11]), .CK(clk), .RN(n770), 
        .Q(work_cntr[11]), .QN(n251) );
  DFFRX2 \write_cntr_reg/q_reg[12]  ( .D(n487), .CK(clk), .RN(n133), .Q(
        write_cntr[12]), .QN(n265) );
  ADDFX2 \DP_OP_229J1_126_7015/U5  ( .A(\DP_OP_229J1_126_7015/n5 ), .B(N89), 
        .CI(\DP_OP_229J1_126_7015/n17 ), .CO(\DP_OP_229J1_126_7015/n4 ), .S(
        N1142) );
  OR2X1 U3 ( .A(work_cntr[13]), .B(n2415), .Y(n2) );
  OR2X1 U4 ( .A(n1812), .B(n2768), .Y(n3) );
  NOR2X1 U5 ( .A(n1704), .B(n1699), .Y(n1710) );
  OR2X1 U6 ( .A(n199), .B(n1567), .Y(n1559) );
  NOR2X1 U7 ( .A(n1726), .B(n1725), .Y(n1734) );
  CLKINVX1 U8 ( .A(next_cr_x[5]), .Y(n1933) );
  OA22X1 U9 ( .A0(n150), .A1(n1), .B0(n151), .B1(n2406), .Y(n2420) );
  OA21XL U10 ( .A0(work_cntr[15]), .A1(n2421), .B0(n2405), .Y(n1) );
  OAI2BB1X1 U11 ( .A0N(n2), .A1N(work_cntr[14]), .B0(n2393), .Y(n2421) );
  NAND3X1 U12 ( .A(write_addr[12]), .B(write_addr[11]), .C(n2848), .Y(n2820)
         );
  OAI31X1 U13 ( .A0(n1868), .A1(n1885), .A2(n1890), .B0(n1887), .Y(n1889) );
  NAND2X1 U14 ( .A(n2272), .B(n2271), .Y(n2264) );
  NOR2BX1 U15 ( .AN(n2200), .B(n2201), .Y(n2222) );
  OAI2BB1X1 U16 ( .A0N(n289), .A1N(n1915), .B0(n2837), .Y(n2835) );
  NOR2X1 U17 ( .A(n229), .B(n255), .Y(n789) );
  OAI2BB1X1 U18 ( .A0N(n3), .A1N(n280), .B0(n1815), .Y(n2775) );
  NOR2BX1 U19 ( .AN(n2290), .B(next_work_cntr[3]), .Y(n2306) );
  OR2X4 U20 ( .A(\DP_OP_590J1_137_6981/I5 ), .B(si_sel), .Y(n729) );
  NOR2X1 U21 ( .A(n1645), .B(n1401), .Y(n1643) );
  NAND2X1 U22 ( .A(n320), .B(global_cntr[5]), .Y(n782) );
  NOR2X1 U23 ( .A(n782), .B(n244), .Y(n326) );
  NOR2X1 U24 ( .A(n319), .B(n242), .Y(n320) );
  BUFX4 U25 ( .A(n2785), .Y(n135) );
  NOR2X1 U26 ( .A(n1774), .B(n318), .Y(expand_sel[2]) );
  OR2X2 U27 ( .A(n789), .B(n748), .Y(en_so) );
  OR2X1 U28 ( .A(n5), .B(n318), .Y(n4) );
  OR2X1 U29 ( .A(n7), .B(n318), .Y(n6) );
  OR2X1 U30 ( .A(n303), .B(n318), .Y(n8) );
  OR2X1 U31 ( .A(n10), .B(n318), .Y(n9) );
  XNOR2X1 U32 ( .A(\DP_OP_229J1_126_7015/n1 ), .B(\DP_OP_229J1_126_7015/n21 ), 
        .Y(n10) );
  AOI21X1 U33 ( .A0(n729), .A1(\C159/DATA3_0 ), .B0(n12), .Y(\im_a[0]_BAR ) );
  AO22X1 U34 ( .A0(n311), .A1(N1347), .B0(n746), .B1(global_cntr[0]), .Y(n12)
         );
  AOI21X1 U35 ( .A0(n729), .A1(\C159/DATA3_1 ), .B0(n14), .Y(\im_a[1]_BAR ) );
  AO22X1 U36 ( .A0(n311), .A1(N1348), .B0(n746), .B1(global_cntr[1]), .Y(n14)
         );
  AOI21X1 U37 ( .A0(n729), .A1(\C159/DATA3_2 ), .B0(n16), .Y(\im_a[2]_BAR ) );
  AO22X1 U38 ( .A0(n728), .A1(N1349), .B0(n746), .B1(global_cntr[2]), .Y(n16)
         );
  AOI21X1 U39 ( .A0(n729), .A1(\C159/DATA3_3 ), .B0(n19), .Y(\im_a[3]_BAR ) );
  AO22X1 U40 ( .A0(n311), .A1(N1350), .B0(n746), .B1(global_cntr[3]), .Y(n19)
         );
  AOI21X1 U41 ( .A0(n729), .A1(\C159/DATA3_4 ), .B0(n21), .Y(\im_a[4]_BAR ) );
  AO22X1 U42 ( .A0(n728), .A1(N1351), .B0(n746), .B1(global_cntr[4]), .Y(n21)
         );
  AOI21X1 U43 ( .A0(n729), .A1(\C159/DATA3_5 ), .B0(n23), .Y(\im_a[5]_BAR ) );
  AO22X1 U44 ( .A0(n311), .A1(N1352), .B0(n746), .B1(global_cntr[5]), .Y(n23)
         );
  AOI21X1 U45 ( .A0(n729), .A1(\C159/DATA3_6 ), .B0(n25), .Y(\im_a[6]_BAR ) );
  AO22X1 U46 ( .A0(n728), .A1(N1353), .B0(n746), .B1(global_cntr[6]), .Y(n25)
         );
  AOI21X1 U47 ( .A0(n729), .A1(\C159/DATA3_7 ), .B0(n29), .Y(\im_a[7]_BAR ) );
  AO22X1 U48 ( .A0(n311), .A1(N1354), .B0(n746), .B1(global_cntr[7]), .Y(n29)
         );
  AOI21X1 U49 ( .A0(n729), .A1(\C159/DATA3_8 ), .B0(n31), .Y(\im_a[8]_BAR ) );
  AO22X1 U50 ( .A0(n728), .A1(N1355), .B0(n746), .B1(global_cntr[8]), .Y(n31)
         );
  AOI21X1 U51 ( .A0(n729), .A1(\C159/DATA3_9 ), .B0(n33), .Y(\im_a[9]_BAR ) );
  AO22X1 U52 ( .A0(n311), .A1(N1356), .B0(n746), .B1(global_cntr[9]), .Y(n33)
         );
  AOI21X1 U53 ( .A0(n729), .A1(\C159/DATA3_10 ), .B0(n35), .Y(\im_a[10]_BAR )
         );
  AO22X1 U54 ( .A0(n728), .A1(N1357), .B0(n746), .B1(global_cntr[10]), .Y(n35)
         );
  AOI21X1 U55 ( .A0(n729), .A1(\C159/DATA3_11 ), .B0(n37), .Y(\im_a[11]_BAR )
         );
  AO22X1 U56 ( .A0(n311), .A1(N1358), .B0(n746), .B1(global_cntr[11]), .Y(n37)
         );
  AOI21X1 U57 ( .A0(n729), .A1(\C159/DATA3_12 ), .B0(n39), .Y(\im_a[12]_BAR )
         );
  AO22X1 U58 ( .A0(n728), .A1(N1359), .B0(n746), .B1(global_cntr[12]), .Y(n39)
         );
  AOI21X1 U59 ( .A0(n729), .A1(\C159/DATA3_13 ), .B0(n41), .Y(\im_a[13]_BAR )
         );
  AO22X1 U60 ( .A0(n311), .A1(N1360), .B0(n746), .B1(global_cntr[13]), .Y(n41)
         );
  AOI21X1 U61 ( .A0(n729), .A1(\C159/DATA3_14 ), .B0(n43), .Y(\im_a[14]_BAR )
         );
  AO22X1 U62 ( .A0(n728), .A1(N1361), .B0(n746), .B1(global_cntr[14]), .Y(n43)
         );
  AOI21X1 U63 ( .A0(n729), .A1(\C159/DATA3_15 ), .B0(n45), .Y(\im_a[15]_BAR )
         );
  AO22X1 U64 ( .A0(n311), .A1(N1362), .B0(n746), .B1(global_cntr[15]), .Y(n45)
         );
  AOI21X1 U65 ( .A0(n729), .A1(\C159/DATA3_16 ), .B0(n47), .Y(\im_a[16]_BAR )
         );
  AO22X1 U66 ( .A0(n728), .A1(N1363), .B0(n746), .B1(global_cntr[16]), .Y(n47)
         );
  AOI21X1 U67 ( .A0(n729), .A1(\C159/DATA3_17 ), .B0(n49), .Y(\im_a[17]_BAR )
         );
  AO22X1 U68 ( .A0(n311), .A1(N1364), .B0(n746), .B1(global_cntr[17]), .Y(n49)
         );
  AOI21X1 U69 ( .A0(n729), .A1(\C159/DATA3_18 ), .B0(n51), .Y(\im_a[18]_BAR )
         );
  AO22X1 U70 ( .A0(n728), .A1(N1365), .B0(n746), .B1(global_cntr[18]), .Y(n51)
         );
  CLKINVX1 U71 ( .A(n2658), .Y(n138) );
  INVX4 U72 ( .A(si_sel), .Y(n318) );
  AND2X2 U73 ( .A(n258), .B(en_so), .Y(si_sel) );
  OAI21XL U74 ( .A0(n134), .A1(n2845), .B0(n362), .Y(n476) );
  CLKINVX1 U75 ( .A(n2120), .Y(n136) );
  CLKINVX1 U76 ( .A(n842), .Y(n53) );
  OA21XL U77 ( .A0(n226), .A1(n53), .B0(n843), .Y(n241) );
  AO22X1 U78 ( .A0(n54), .A1(n136), .B0(n2165), .B1(n2120), .Y(n2181) );
  CLKINVX1 U79 ( .A(n2165), .Y(n54) );
  CLKINVX1 U80 ( .A(curr_time[23]), .Y(n55) );
  OAI211X1 U81 ( .A0(curr_time[21]), .A1(n55), .B0(n430), .C0(curr_time[22]), 
        .Y(n56) );
  NAND2X1 U82 ( .A(n431), .B(n56), .Y(n426) );
  NAND2BX1 U83 ( .AN(n1797), .B(n424), .Y(n549) );
  NOR2X1 U84 ( .A(n2832), .B(n282), .Y(n57) );
  OAI21XL U85 ( .A0(write_addr[19]), .A1(n2833), .B0(n740), .Y(n58) );
  NOR2X1 U86 ( .A(n299), .B(n704), .Y(n59) );
  AOI2BB2X1 U87 ( .B0(n159), .B1(n697), .A0N(n718), .A1N(n283), .Y(n60) );
  OAI21XL U88 ( .A0(n710), .A1(n607), .B0(n60), .Y(n61) );
  AOI211X1 U89 ( .A0(n582), .A1(n723), .B0(n59), .C0(n61), .Y(n62) );
  NAND2X1 U90 ( .A(n720), .B(\C158/DATA2_17 ), .Y(n63) );
  OAI211X1 U91 ( .A0(n57), .A1(n58), .B0(n62), .C0(n63), .Y(n64) );
  AO22X1 U92 ( .A0(n314), .A1(n64), .B0(global_cntr[17]), .B1(n724), .Y(
        \C2/Z_17 ) );
  OAI2BB1X1 U93 ( .A0N(n853), .A1N(n241), .B0(n857), .Y(n2720) );
  NAND2BX1 U94 ( .AN(n1974), .B(n1970), .Y(n1963) );
  OAI211XL U95 ( .A0(n398), .A1(curr_time[10]), .B0(n401), .C0(curr_time[9]), 
        .Y(n65) );
  AND2X1 U96 ( .A(n533), .B(n65), .Y(n539) );
  NAND3X1 U97 ( .A(n548), .B(n547), .C(n549), .Y(n66) );
  NOR2X1 U98 ( .A(n546), .B(n66), .Y(\DP_OP_229J1_126_7015/I2 ) );
  OAI22XL U99 ( .A0(\sftr_n[0]_BAR ), .A1(n223), .B0(n2854), .B1(n651), .Y(n67) );
  AOI22X1 U100 ( .A0(\C158/DATA2_9 ), .A1(n720), .B0(n2856), .B1(n67), .Y(n68)
         );
  OA22X1 U101 ( .A0(n718), .A1(n294), .B0(n719), .B1(n237), .Y(n69) );
  OAI211X1 U102 ( .A0(n650), .A1(n715), .B0(n68), .C0(n69), .Y(n70) );
  AOI21X1 U103 ( .A0(n2858), .A1(n723), .B0(n70), .Y(n71) );
  OAI22XL U104 ( .A0(n1783), .A1(n240), .B0(n725), .B1(n71), .Y(\C2/Z_9 ) );
  OAI21XL U105 ( .A0(n2782), .A1(n2784), .B0(n744), .Y(n72) );
  AOI21X1 U106 ( .A0(n2784), .A1(write_addr[19]), .B0(n72), .Y(n582) );
  OAI2BB1X1 U107 ( .A0N(n2545), .A1N(n141), .B0(n2542), .Y(n2543) );
  AO22X1 U108 ( .A0(n2722), .A1(n73), .B0(n2724), .B1(n233), .Y(n2727) );
  CLKINVX1 U109 ( .A(n2723), .Y(n73) );
  AOI2BB1X1 U110 ( .A0N(write_cntr[12]), .A1N(n1560), .B0(n279), .Y(n1573) );
  OAI211X1 U111 ( .A0(n1734), .A1(n212), .B0(n1732), .C0(n1729), .Y(n74) );
  AOI31X1 U112 ( .A0(n1728), .A1(n1731), .A2(n74), .B0(n1727), .Y(n1733) );
  NOR2XL U113 ( .A(n2121), .B(n2159), .Y(n75) );
  AOI31X1 U114 ( .A0(n2118), .A1(n2191), .A2(n75), .B0(n2134), .Y(n2133) );
  OAI2BB1X1 U115 ( .A0N(n456), .A1N(n457), .B0(n458), .Y(n460) );
  NOR4X1 U116 ( .A(global_cntr[9]), .B(global_cntr[16]), .C(global_cntr[14]), 
        .D(global_cntr[17]), .Y(n76) );
  NOR4X1 U117 ( .A(global_cntr[3]), .B(global_cntr[5]), .C(global_cntr[6]), 
        .D(global_cntr[4]), .Y(n77) );
  NAND3X1 U118 ( .A(n1553), .B(n76), .C(n77), .Y(n78) );
  NOR3X1 U119 ( .A(global_cntr[19]), .B(global_cntr[18]), .C(n78), .Y(n1554)
         );
  AO21X1 U120 ( .A0(\DP_OP_229J1_126_7015/n24 ), .A1(n173), .B0(
        \DP_OP_229J1_126_7015/I2 ), .Y(n79) );
  AND2X1 U121 ( .A(\DP_OP_229J1_126_7015/n4 ), .B(n79), .Y(
        \DP_OP_229J1_126_7015/n3 ) );
  AOI2BB2X1 U122 ( .B0(\DP_OP_229J1_126_7015/n4 ), .B1(n79), .A0N(
        \DP_OP_229J1_126_7015/n4 ), .A1N(n79), .Y(N1143) );
  OA22X1 U123 ( .A0(n718), .A1(n236), .B0(n719), .B1(n2811), .Y(n80) );
  NAND2X1 U124 ( .A(write_addr[1]), .B(n720), .Y(n81) );
  OAI211X1 U125 ( .A0(n717), .A1(write_addr[1]), .B0(n80), .C0(n81), .Y(n82)
         );
  OAI22XL U126 ( .A0(n288), .A1(n721), .B0(n716), .B1(n715), .Y(n83) );
  AOI211X1 U127 ( .A0(n723), .A1(n722), .B0(n82), .C0(n83), .Y(n84) );
  OAI22XL U128 ( .A0(n253), .A1(n1783), .B0(n313), .B1(n84), .Y(n85) );
  AOI22X1 U129 ( .A0(N1347), .A1(n312), .B0(\DP_OP_590J1_137_6981/I5 ), .B1(
        n85), .Y(n86) );
  NAND2BX1 U130 ( .AN(n313), .B(curr_photo_addr[0]), .Y(n87) );
  NOR2X1 U131 ( .A(n86), .B(n87), .Y(\DP_OP_590J1_137_6981/n20 ) );
  AOI2BB2X1 U132 ( .B0(n86), .B1(n87), .A0N(n86), .A1N(n87), .Y(\C159/DATA3_0 ) );
  OAI2BB2XL U133 ( .B0(n741), .B1(n2785), .A0N(n135), .A1N(n690), .Y(n478) );
  INVXL U134 ( .A(n2546), .Y(n88) );
  CLKINVX1 U135 ( .A(n141), .Y(n89) );
  AOI32X1 U136 ( .A0(n2545), .A1(n141), .A2(n88), .B0(n2547), .B1(n89), .Y(
        n2554) );
  OAI2BB1X1 U137 ( .A0N(n196), .A1N(n1694), .B0(n1686), .Y(n90) );
  AOI2BB2X1 U138 ( .B0(n1687), .B1(n90), .A0N(n1687), .A1N(n90), .Y(n1690) );
  OAI2BB1X1 U139 ( .A0N(n2581), .A1N(n2586), .B0(n2578), .Y(n2579) );
  AOI2BB2X1 U140 ( .B0(n153), .B1(n137), .A0N(n153), .A1N(n137), .Y(n91) );
  OAI2BB1X1 U141 ( .A0N(n1719), .A1N(n1712), .B0(n1720), .Y(n92) );
  CLKINVX1 U142 ( .A(n1712), .Y(n93) );
  AOI31X1 U143 ( .A0(n1721), .A1(n91), .A2(n92), .B0(n93), .Y(n1715) );
  NOR2X1 U144 ( .A(n1982), .B(n1992), .Y(n94) );
  NAND2X1 U145 ( .A(n1978), .B(n94), .Y(n1983) );
  AOI21X1 U146 ( .A0(n2728), .A1(n2726), .B0(n2732), .Y(n2734) );
  AOI21X1 U147 ( .A0(n1596), .A1(n1603), .B0(n95), .Y(n1594) );
  CLKINVX1 U148 ( .A(n1601), .Y(n95) );
  OAI2BB1X1 U149 ( .A0N(n350), .A1N(\s_1[3] ), .B0(n986), .Y(n411) );
  NAND2X1 U150 ( .A(n1745), .B(n1735), .Y(n96) );
  NOR2X1 U151 ( .A(n1738), .B(n96), .Y(n1739) );
  NOR2X1 U152 ( .A(n2744), .B(n1873), .Y(n97) );
  XNOR2X1 U153 ( .A(n97), .B(n913), .Y(n927) );
  AOI31X1 U154 ( .A0(n826), .A1(next_cr_x[6]), .A2(n824), .B0(n823), .Y(n1021)
         );
  OAI2BB1X1 U155 ( .A0N(n2196), .A1N(n2199), .B0(n2198), .Y(n2180) );
  OAI2BB1X1 U156 ( .A0N(n342), .A1N(m_1[3]), .B0(n979), .Y(n394) );
  NOR4BX1 U157 ( .AN(n142), .B(n2217), .C(n2237), .D(n2232), .Y(n98) );
  NAND4BX1 U158 ( .AN(n2245), .B(n98), .C(n2259), .D(n2248), .Y(n2246) );
  OAI2BB1X1 U159 ( .A0N(n2031), .A1N(n2030), .B0(n2032), .Y(n99) );
  XNOR2X1 U160 ( .A(n99), .B(n2033), .Y(n2034) );
  OAI2BB1X1 U161 ( .A0N(n2619), .A1N(n2624), .B0(n2616), .Y(n2617) );
  AOI2BB1X1 U162 ( .A0N(n1813), .A1N(n282), .B0(n2855), .Y(n1823) );
  NAND3X1 U163 ( .A(n2334), .B(n2307), .C(n2308), .Y(n2314) );
  AO21X1 U164 ( .A0(\DP_OP_229J1_126_7015/n25 ), .A1(n173), .B0(
        \DP_OP_229J1_126_7015/I2 ), .Y(n100) );
  AND2X1 U165 ( .A(\DP_OP_229J1_126_7015/n3 ), .B(n100), .Y(
        \DP_OP_229J1_126_7015/n2 ) );
  AOI2BB2X1 U166 ( .B0(\DP_OP_229J1_126_7015/n3 ), .B1(n100), .A0N(
        \DP_OP_229J1_126_7015/n3 ), .A1N(n100), .Y(N1144) );
  NOR3XL U167 ( .A(n754), .B(n755), .C(n756), .Y(n101) );
  NOR3X1 U168 ( .A(n753), .B(n751), .C(n752), .Y(n102) );
  NAND4X1 U169 ( .A(n795), .B(n784), .C(n101), .D(n102), .Y(n785) );
  NOR2BX1 U170 ( .AN(n742), .B(n2867), .Y(n737) );
  OAI2BB2XL U171 ( .B0(n2785), .B1(n223), .A0N(n2858), .A1N(n135), .Y(n442) );
  OAI2BB1X1 U172 ( .A0N(n2526), .A1N(n2531), .B0(n2523), .Y(n2524) );
  OAI2BB1X1 U173 ( .A0N(n2562), .A1N(n2567), .B0(n149), .Y(n2560) );
  NAND2X1 U174 ( .A(n1962), .B(n1970), .Y(n103) );
  OAI21XL U175 ( .A0(n1982), .A1(n1981), .B0(n1964), .Y(n104) );
  XNOR2X1 U176 ( .A(n104), .B(n103), .Y(n1979) );
  NAND3BX1 U177 ( .AN(n907), .B(n902), .C(n905), .Y(n903) );
  CLKINVX1 U178 ( .A(n2726), .Y(n105) );
  AOI32X1 U179 ( .A0(n2728), .A1(n105), .A2(n2727), .B0(n2726), .B1(n2725), 
        .Y(n2731) );
  OAI2BB1X1 U180 ( .A0N(n1572), .A1N(n1573), .B0(n1563), .Y(n1621) );
  AOI2BB1X1 U181 ( .A0N(n1738), .A1N(n1737), .B0(n1734), .Y(n106) );
  NAND2X1 U182 ( .A(n1731), .B(n1732), .Y(n107) );
  AOI2BB2X1 U183 ( .B0(n106), .B1(n107), .A0N(n106), .A1N(n107), .Y(n1736) );
  OAI2BB1X1 U184 ( .A0N(n2600), .A1N(n2605), .B0(n2597), .Y(n2598) );
  CLKINVX1 U185 ( .A(curr_time[4]), .Y(n108) );
  NAND2X1 U186 ( .A(n353), .B(n411), .Y(n109) );
  OAI211X1 U187 ( .A0(n986), .A1(n108), .B0(n989), .C0(n109), .Y(n413) );
  OAI2BB1X1 U188 ( .A0N(n1617), .A1N(n1618), .B0(n155), .Y(n1798) );
  NAND3BX1 U189 ( .AN(n829), .B(n1018), .C(n1015), .Y(n824) );
  NOR2X1 U190 ( .A(n2190), .B(n2177), .Y(n110) );
  OAI2BB2XL U191 ( .B0(n2176), .B1(n110), .A0N(n2211), .A1N(n2212), .Y(n111)
         );
  NAND2X1 U192 ( .A(n2207), .B(n111), .Y(n2215) );
  OAI2BB1X1 U193 ( .A0N(n427), .A1N(n426), .B0(n973), .Y(n456) );
  CLKINVX1 U194 ( .A(curr_time[12]), .Y(n112) );
  NAND2X1 U195 ( .A(n345), .B(n394), .Y(n113) );
  OAI211X1 U196 ( .A0(n979), .A1(n112), .B0(n982), .C0(n113), .Y(n392) );
  NAND2BX1 U197 ( .AN(n717), .B(n2847), .Y(n651) );
  OAI21XL U198 ( .A0(n1932), .A1(n1866), .B0(n1865), .Y(n114) );
  NAND2X1 U199 ( .A(n1867), .B(n114), .Y(n1890) );
  AOI2BB2X1 U200 ( .B0(write_addr[19]), .B1(fb_addr[19]), .A0N(write_addr[19]), 
        .A1N(fb_addr[19]), .Y(n115) );
  AOI2BB2X1 U201 ( .B0(\DP_OP_590J1_137_6981/n22 ), .B1(n115), .A0N(
        \DP_OP_590J1_137_6981/n22 ), .A1N(n115), .Y(N1366) );
  OAI2BB1X1 U202 ( .A0N(n1278), .A1N(n1262), .B0(n1267), .Y(n116) );
  NAND2X1 U203 ( .A(n1279), .B(n116), .Y(n117) );
  OAI211X1 U204 ( .A0(n1279), .A1(n116), .B0(n1557), .C0(n117), .Y(n384) );
  AO21X1 U205 ( .A0(n118), .A1(n2837), .B0(n2836), .Y(n683) );
  CLKINVX1 U206 ( .A(write_addr[4]), .Y(n118) );
  OAI21XL U207 ( .A0(n2260), .A1(n2221), .B0(n2226), .Y(n119) );
  XNOR2X1 U208 ( .A(n119), .B(n2222), .Y(n2289) );
  OA21XL U209 ( .A0(n2451), .A1(n2450), .B0(n2449), .Y(n120) );
  AOI2BB1X1 U210 ( .A0N(work_cntr[9]), .A1N(n2462), .B0(n2452), .Y(n121) );
  AOI2BB2X1 U211 ( .B0(n120), .B1(n121), .A0N(n120), .A1N(n2453), .Y(n2463) );
  OAI21XL U212 ( .A0(n2060), .A1(n2059), .B0(n2063), .Y(n122) );
  NAND3X1 U213 ( .A(n2065), .B(n2057), .C(n122), .Y(n123) );
  AOI32X1 U214 ( .A0(n2065), .A1(n123), .A2(n2054), .B0(n2058), .B1(n123), .Y(
        n2061) );
  AOI21X1 U215 ( .A0(n2267), .A1(n2291), .B0(n211), .Y(n210) );
  AO21X1 U216 ( .A0(\DP_OP_229J1_126_7015/n26 ), .A1(n173), .B0(
        \DP_OP_229J1_126_7015/I2 ), .Y(n124) );
  AND2X1 U217 ( .A(\DP_OP_229J1_126_7015/n2 ), .B(n124), .Y(
        \DP_OP_229J1_126_7015/n1 ) );
  AOI2BB2X1 U218 ( .B0(\DP_OP_229J1_126_7015/n2 ), .B1(n124), .A0N(
        \DP_OP_229J1_126_7015/n2 ), .A1N(n124), .Y(N1145) );
  NOR2X1 U219 ( .A(n2306), .B(n2308), .Y(n125) );
  AOI2BB2X1 U220 ( .B0(n2307), .B1(n125), .A0N(n2307), .A1N(n125), .Y(n2333)
         );
  OAI2BB1X1 U221 ( .A0N(n2636), .A1N(n2641), .B0(n2635), .Y(n2645) );
  OAI21XL U222 ( .A0(n1676), .A1(n1677), .B0(n1670), .Y(n126) );
  NAND2X1 U223 ( .A(n1669), .B(n126), .Y(n1686) );
  NAND2X1 U224 ( .A(n303), .B(n2695), .Y(n127) );
  OAI22XL U225 ( .A0(n2686), .A1(n127), .B0(n2685), .B1(n303), .Y(n452) );
  AOI21X1 U226 ( .A0(n305), .A1(n2793), .B0(n2792), .Y(next_photo[0]) );
  CLKINVX1 U227 ( .A(n801), .Y(n128) );
  OAI211X1 U228 ( .A0(n1783), .A1(n128), .B0(n802), .C0(n1787), .Y(
        next_state[1]) );
  NOR2BX1 U229 ( .AN(n781), .B(n782), .Y(n129) );
  AOI2BB1X1 U230 ( .A0N(global_cntr[6]), .A1N(n129), .B0(n326), .Y(n756) );
  OAI2BB2XL U231 ( .B0(n2785), .B1(n296), .A0N(n2828), .A1N(n135), .Y(n440) );
  NOR3X2 U232 ( .A(n2124), .B(n2112), .C(n2115), .Y(n130) );
  OR2X1 U233 ( .A(n215), .B(n1856), .Y(n131) );
  CLKINVX1 U234 ( .A(n2011), .Y(n167) );
  OAI21X1 U235 ( .A0(n1458), .A1(n1462), .B0(n1457), .Y(n132) );
  NAND2BX1 U236 ( .AN(n2381), .B(n2417), .Y(n2415) );
  NOR2X1 U237 ( .A(n1857), .B(n1941), .Y(n1856) );
  OA21X2 U238 ( .A0(n251), .A1(n1455), .B0(n1450), .Y(n1458) );
  AOI32X1 U239 ( .A0(n1768), .A1(n1788), .A2(n232), .B0(n1776), .B1(n1788), 
        .Y(n1790) );
  NOR2X1 U240 ( .A(n1005), .B(n266), .Y(n1004) );
  OAI22X2 U241 ( .A0(n1804), .A1(n2725), .B0(n877), .B1(n2728), .Y(n894) );
  OAI22X2 U242 ( .A0(write_cntr[8]), .A1(n830), .B0(n269), .B1(n838), .Y(n877)
         );
  NAND2X1 U243 ( .A(n1772), .B(n263), .Y(n1780) );
  NOR2X2 U244 ( .A(n2291), .B(n2267), .Y(n211) );
  NAND2X2 U245 ( .A(n1643), .B(n259), .Y(n1788) );
  BUFX4 U246 ( .A(n770), .Y(n133) );
  INVX12 U247 ( .A(reset), .Y(n770) );
  OAI31X1 U248 ( .A0(n1745), .A1(n1744), .A2(n1743), .B0(n1742), .Y(n1749) );
  INVX6 U249 ( .A(n135), .Y(n134) );
  NAND2X4 U250 ( .A(n313), .B(n1783), .Y(\DP_OP_590J1_137_6981/I5 ) );
  AOI221X1 U251 ( .A0(n2289), .A1(n2288), .B0(n2287), .B1(n2288), .C0(n2295), 
        .Y(n2317) );
  NOR2X1 U252 ( .A(n2077), .B(n2076), .Y(n2089) );
  NOR2X1 U253 ( .A(n142), .B(n2223), .Y(n2261) );
  OAI21X1 U254 ( .A0(n2748), .A1(n2747), .B0(n2746), .Y(n2753) );
  OR2XL U255 ( .A(n193), .B(n138), .Y(n192) );
  OAI21X1 U256 ( .A0(n2654), .A1(n2653), .B0(n2652), .Y(n2660) );
  OAI21X1 U257 ( .A0(n2730), .A1(n2731), .B0(n2729), .Y(n2738) );
  NOR2X1 U258 ( .A(n1859), .B(n1846), .Y(n1847) );
  OAI21X1 U259 ( .A0(n872), .A1(n871), .B0(n870), .Y(n883) );
  OAI21X1 U260 ( .A0(n266), .A1(n1478), .B0(n1477), .Y(n1484) );
  NOR2X1 U261 ( .A(n268), .B(n1092), .Y(n1110) );
  OAI21X1 U262 ( .A0(n2452), .A1(n2453), .B0(n2457), .Y(n2456) );
  NAND2X1 U263 ( .A(n316), .B(n2552), .Y(n2116) );
  NAND2X1 U264 ( .A(n316), .B(n2637), .Y(n2265) );
  NAND2X1 U265 ( .A(n316), .B(n2571), .Y(n2145) );
  NOR2X2 U266 ( .A(n317), .B(n2581), .Y(next_work_cntr[10]) );
  OAI21X1 U267 ( .A0(n1282), .A1(n257), .B0(n1284), .Y(n1299) );
  OAI22X1 U268 ( .A0(n2433), .A1(work_cntr[10]), .B0(n2432), .B1(n228), .Y(
        n2450) );
  NOR2X1 U269 ( .A(n1401), .B(n1284), .Y(n1292) );
  OAI22X1 U270 ( .A0(n1355), .A1(n268), .B0(n1354), .B1(n1723), .Y(n1372) );
  NOR2X1 U271 ( .A(n1818), .B(n222), .Y(n1817) );
  NAND2X1 U272 ( .A(curr_time[15]), .B(n978), .Y(n345) );
  NAND2X1 U273 ( .A(curr_time[7]), .B(n985), .Y(n353) );
  NOR2X2 U274 ( .A(\state[2] ), .B(n26), .Y(n748) );
  AOI211X1 U275 ( .A0(n744), .A1(n2681), .B0(n310), .C0(n2683), .Y(n2876) );
  OA21XL U276 ( .A0(n1913), .A1(n1926), .B0(n1912), .Y(n1923) );
  AOI221X1 U277 ( .A0(n1908), .A1(n1907), .B0(n1906), .B1(n1907), .C0(n1920), 
        .Y(n1909) );
  AND2X2 U278 ( .A(n1906), .B(n1919), .Y(\next_cr_y[0] ) );
  NAND2X2 U279 ( .A(im_wen_n), .B(n316), .Y(n2785) );
  OAI31X1 U280 ( .A0(n959), .A1(n966), .A2(n963), .B0(n958), .Y(n1906) );
  OAI2BB2X1 U281 ( .B0(n1222), .B1(n1211), .A0N(n1222), .A1N(n1211), .Y(n1250)
         );
  NOR2X1 U282 ( .A(n271), .B(n2794), .Y(n1796) );
  OA21XL U283 ( .A0(n2641), .A1(n2640), .B0(n2639), .Y(n2650) );
  OAI31X1 U284 ( .A0(n1531), .A1(N1826), .A2(n1530), .B0(n1529), .Y(n1537) );
  OA21XL U285 ( .A0(n2624), .A1(n2623), .B0(n2622), .Y(n2630) );
  OA21XL U286 ( .A0(n1504), .A1(n1503), .B0(n1502), .Y(n1511) );
  OA21XL U287 ( .A0(n1979), .A1(n1978), .B0(n1980), .Y(n2000) );
  OAI31X1 U288 ( .A0(n860), .A1(n859), .A2(n2719), .B0(n858), .Y(n872) );
  OAI31X1 U289 ( .A0(n1493), .A1(work_cntr[6]), .A2(n1492), .B0(n1491), .Y(
        n1498) );
  OAI211X1 U290 ( .A0(n1956), .A1(n1744), .B0(n1748), .C0(n1745), .Y(n1742) );
  AND4X1 U291 ( .A(n556), .B(n555), .C(n554), .D(n553), .Y(
        \DP_OP_229J1_126_7015/I3 ) );
  OA21XL U292 ( .A0(n2586), .A1(n2585), .B0(n2584), .Y(n2592) );
  OAI211X1 U293 ( .A0(n1972), .A1(n1961), .B0(n1962), .C0(n1971), .Y(n1964) );
  OAI211X1 U294 ( .A0(n1708), .A1(n1716), .B0(n1712), .C0(n1719), .Y(n1728) );
  OAI21XL U295 ( .A0(n261), .A1(n1470), .B0(n1465), .Y(n1473) );
  OAI31X1 U296 ( .A0(n1096), .A1(n1095), .A2(n1094), .B0(n1093), .Y(n1136) );
  AND2XL U297 ( .A(n316), .B(n2628), .Y(n2224) );
  CLKINVX1 U298 ( .A(n1710), .Y(n137) );
  AOI22X1 U299 ( .A0(\state[2] ), .A1(n799), .B0(n807), .B1(n803), .Y(n2086)
         );
  NAND2X1 U300 ( .A(n258), .B(n804), .Y(n807) );
  OAI21XL U301 ( .A0(n2539), .A1(n2540), .B0(n2538), .Y(n2548) );
  OA21XL U302 ( .A0(n1442), .A1(n1446), .B0(n1441), .Y(n1448) );
  OR2XL U303 ( .A(n757), .B(n785), .Y(n195) );
  OR2XL U304 ( .A(n750), .B(n749), .Y(n194) );
  AOI31X1 U305 ( .A0(curr_time[1]), .A1(n417), .A2(n191), .B0(n524), .Y(n545)
         );
  OR2X1 U306 ( .A(n200), .B(n201), .Y(n197) );
  AOI211X1 U307 ( .A0(n1292), .A1(work_cntr[19]), .B0(n1287), .C0(n1286), .Y(
        n1297) );
  AOI211X1 U308 ( .A0(n1032), .A1(n1033), .B0(n561), .C0(n558), .Y(n562) );
  XOR2X1 U309 ( .A(n426), .B(curr_time[20]), .Y(n976) );
  OA21XL U310 ( .A0(n2460), .A1(n221), .B0(n2459), .Y(n2482) );
  OR2X1 U311 ( .A(n213), .B(n214), .Y(n212) );
  NAND2BX4 U312 ( .AN(n27), .B(n338), .Y(n1783) );
  NOR2X1 U313 ( .A(\state[2] ), .B(n255), .Y(n338) );
  INVX1 U314 ( .A(curr_photo_size[0]), .Y(n378) );
  INVX1 U315 ( .A(curr_photo_size[1]), .Y(n775) );
  CLKINVX1 U316 ( .A(n1473), .Y(n140) );
  CLKINVX1 U317 ( .A(n2548), .Y(n141) );
  NAND2X1 U318 ( .A(n2371), .B(n2372), .Y(n2330) );
  OAI31X1 U319 ( .A0(n886), .A1(n885), .A2(n2725), .B0(n884), .Y(n897) );
  AND2X2 U320 ( .A(n874), .B(n1804), .Y(n886) );
  CLKINVX1 U321 ( .A(n2224), .Y(n142) );
  NAND2X1 U322 ( .A(n843), .B(n842), .Y(n849) );
  CLKINVX1 U323 ( .A(n841), .Y(n843) );
  NAND2X2 U324 ( .A(n231), .B(n252), .Y(n1401) );
  NAND2BX1 U325 ( .AN(n1210), .B(n1203), .Y(n1220) );
  NOR2X1 U326 ( .A(n1574), .B(n1576), .Y(n1583) );
  NAND2X1 U327 ( .A(n2383), .B(n1328), .Y(n1284) );
  NOR2X1 U328 ( .A(n1354), .B(n1709), .Y(n1328) );
  NAND2BX1 U329 ( .AN(n1252), .B(n1238), .Y(n1246) );
  OAI2BB2X1 U330 ( .B0(n1235), .B1(n1234), .A0N(n1235), .A1N(n1234), .Y(n1252)
         );
  CLKINVX1 U331 ( .A(n2378), .Y(n2496) );
  OAI21X1 U332 ( .A0(n270), .A1(n1514), .B0(n1513), .Y(n1517) );
  OAI21X1 U333 ( .A0(n2636), .A1(n2644), .B0(n2640), .Y(n2642) );
  OAI21X1 U334 ( .A0(n221), .A1(n1506), .B0(n1503), .Y(n1500) );
  NAND4X1 U335 ( .A(N1139), .B(N1138), .C(N1140), .D(cr_read_cntr[3]), .Y(
        n2689) );
  OAI21X1 U336 ( .A0(n1137), .A1(n1136), .B0(n1135), .Y(n1144) );
  OAI21X1 U337 ( .A0(n2475), .A1(n2483), .B0(n164), .Y(n2478) );
  OAI211X1 U338 ( .A0(n2385), .A1(work_cntr[19]), .B0(n2388), .C0(n2384), .Y(
        n2389) );
  CLKINVX1 U339 ( .A(n2386), .Y(n2385) );
  OAI21X1 U340 ( .A0(n2567), .A1(n2566), .B0(n2565), .Y(n2573) );
  INVXL U341 ( .A(n2592), .Y(n143) );
  INVXL U342 ( .A(n2650), .Y(n144) );
  OAI21X1 U343 ( .A0(n2605), .A1(n2604), .B0(n2603), .Y(n2611) );
  INVXL U344 ( .A(n2630), .Y(n145) );
  NOR2X1 U345 ( .A(work_cntr[4]), .B(n317), .Y(n2068) );
  INVXL U346 ( .A(n1448), .Y(n146) );
  INVXL U347 ( .A(n1511), .Y(n147) );
  OAI21X1 U348 ( .A0(n2531), .A1(n2530), .B0(n2529), .Y(n2537) );
  NAND2X1 U349 ( .A(n832), .B(n831), .Y(n1019) );
  NAND2X1 U350 ( .A(n832), .B(n822), .Y(n831) );
  OAI21X1 U351 ( .A0(n2395), .A1(n257), .B0(n2394), .Y(n2396) );
  OAI21X1 U352 ( .A0(n2827), .A1(n2853), .B0(n2851), .Y(n2825) );
  OAI21X1 U353 ( .A0(n2301), .A1(n2300), .B0(n2325), .Y(n2323) );
  NAND4BX1 U354 ( .AN(n2315), .B(n2313), .C(n2317), .D(n2293), .Y(n2300) );
  OAI211X1 U355 ( .A0(n988), .A1(n553), .B0(n519), .C0(n518), .Y(\C1/Z_2 ) );
  OAI21X1 U356 ( .A0(n2437), .A1(n2431), .B0(n2441), .Y(n2443) );
  OAI21X1 U357 ( .A0(n905), .A1(n904), .B0(n903), .Y(n910) );
  OAI21X1 U358 ( .A0(n2648), .A1(n2652), .B0(n2647), .Y(n2656) );
  AOI31X1 U359 ( .A0(n1632), .A1(n1624), .A2(n1634), .B0(n1614), .Y(n1623) );
  AOI2BB2X2 U360 ( .B0(n1119), .B1(n1118), .A0N(n1119), .A1N(n1118), .Y(n1182)
         );
  OAI21X1 U361 ( .A0(n2870), .A1(n2869), .B0(n742), .Y(n2875) );
  AOI2BB2X2 U362 ( .B0(n1832), .B1(n1831), .A0N(n1832), .A1N(n1831), .Y(n1845)
         );
  NOR3X1 U363 ( .A(N1826), .B(N1827), .C(n1788), .Y(n2815) );
  OAI31X1 U364 ( .A0(n1084), .A1(n1062), .A2(n1056), .B0(n1089), .Y(n1088) );
  OAI22X1 U365 ( .A0(n1055), .A1(n1054), .B0(n1053), .B1(n1052), .Y(n1089) );
  OAI22X1 U366 ( .A0(n2016), .A1(n2015), .B0(n167), .B1(n2014), .Y(n2020) );
  INVXL U367 ( .A(n2559), .Y(n148) );
  INVXL U368 ( .A(n148), .Y(n149) );
  OAI31X1 U369 ( .A0(n865), .A1(n864), .A2(n866), .B0(n863), .Y(n878) );
  OAI21X1 U370 ( .A0(n1172), .A1(n1171), .B0(n1170), .Y(n1173) );
  CLKINVX1 U371 ( .A(n1189), .Y(n1171) );
  OAI21X1 U372 ( .A0(n1140), .A1(n1170), .B0(n1139), .Y(n1141) );
  OAI21X1 U373 ( .A0(n2201), .A1(n2226), .B0(n2200), .Y(n2202) );
  CLKINVX1 U374 ( .A(n2216), .Y(n2226) );
  OAI21X1 U375 ( .A0(n1077), .A1(n1100), .B0(n1076), .Y(n1078) );
  OAI21X1 U376 ( .A0(n1590), .A1(n1605), .B0(n1589), .Y(n1591) );
  AOI211X1 U377 ( .A0(n1548), .A1(n1547), .B0(curr_photo_size[0]), .C0(n1546), 
        .Y(n1784) );
  INVXL U378 ( .A(n2407), .Y(n150) );
  INVXL U379 ( .A(n150), .Y(n151) );
  AOI2BB2X2 U380 ( .B0(n1125), .B1(n1124), .A0N(n1125), .A1N(n1124), .Y(n1154)
         );
  NAND2BX2 U381 ( .AN(n1109), .B(n1097), .Y(n1125) );
  AOI2BB2X2 U382 ( .B0(n1377), .B1(n1376), .A0N(n1377), .A1N(n1375), .Y(n1385)
         );
  CLKINVX1 U383 ( .A(n1711), .Y(n152) );
  CLKINVX1 U384 ( .A(n152), .Y(n153) );
  NOR2X1 U385 ( .A(n1039), .B(work_cntr[16]), .Y(n2383) );
  NOR2X1 U386 ( .A(n2044), .B(n2041), .Y(n2045) );
  NOR2X1 U387 ( .A(n1674), .B(n1662), .Y(n1687) );
  NAND2X1 U388 ( .A(n1667), .B(n1675), .Y(n1662) );
  NOR2X1 U389 ( .A(n1763), .B(n1762), .Y(n1779) );
  CLKINVX1 U390 ( .A(n1756), .Y(n1763) );
  OAI211X1 U391 ( .A0(n2742), .A1(n2741), .B0(n2740), .C0(n2739), .Y(n2747) );
  OAI2BB2X1 U392 ( .B0(n2423), .B1(n2415), .A0N(n2423), .A1N(n2415), .Y(n2425)
         );
  OAI31X1 U393 ( .A0(n953), .A1(n952), .A2(n2717), .B0(n951), .Y(n963) );
  NOR2BX1 U394 ( .AN(n1803), .B(n944), .Y(n953) );
  OAI21X1 U395 ( .A0(curr_time[7]), .A1(n773), .B0(n984), .Y(n986) );
  OAI2BB2X1 U396 ( .B0(n1848), .B1(n1925), .A0N(n1847), .A1N(n1941), .Y(n1849)
         );
  AND2X2 U397 ( .A(n413), .B(n412), .Y(n419) );
  OAI31X1 U398 ( .A0(n1453), .A1(work_cntr[11]), .A2(n1452), .B0(n1451), .Y(
        n1460) );
  NAND2X1 U399 ( .A(n1445), .B(n1447), .Y(n1453) );
  OAI31X1 U400 ( .A0(n2536), .A1(n2535), .A2(n2534), .B0(n2533), .Y(n2542) );
  NAND2X1 U401 ( .A(n2524), .B(n2525), .Y(n2536) );
  OAI31X1 U402 ( .A0(n2572), .A1(n2571), .A2(n2570), .B0(n2569), .Y(n2578) );
  NAND2X1 U403 ( .A(n2560), .B(n2561), .Y(n2572) );
  OAI31X1 U404 ( .A0(n1468), .A1(work_cntr[9]), .A2(n1467), .B0(n1466), .Y(
        n1475) );
  NAND2X1 U405 ( .A(n1461), .B(n1463), .Y(n1468) );
  NAND2X1 U406 ( .A(n2617), .B(n2618), .Y(n2629) );
  OAI31X1 U407 ( .A0(n2610), .A1(n2609), .A2(n2608), .B0(n2607), .Y(n2616) );
  NAND2X1 U408 ( .A(n2598), .B(n2599), .Y(n2610) );
  OAI31X1 U409 ( .A0(n2591), .A1(n2590), .A2(n2589), .B0(n2588), .Y(n2597) );
  NAND2X1 U410 ( .A(n2579), .B(n2580), .Y(n2591) );
  OAI21X1 U411 ( .A0(n1641), .A1(n1951), .B0(n1771), .Y(n1775) );
  NAND2X1 U412 ( .A(n2654), .B(n2658), .Y(n1951) );
  CLKINVX1 U413 ( .A(n1192), .Y(n1218) );
  NAND2X1 U414 ( .A(n1171), .B(n1188), .Y(n1192) );
  NOR2X1 U415 ( .A(n234), .B(n1561), .Y(n1571) );
  NAND2X1 U416 ( .A(n856), .B(n864), .Y(n871) );
  INVXL U417 ( .A(n1615), .Y(n154) );
  CLKINVX1 U418 ( .A(n154), .Y(n155) );
  CLKINVX1 U419 ( .A(n817), .Y(n821) );
  NAND4X1 U420 ( .A(write_cntr[8]), .B(write_cntr[7]), .C(write_cntr[6]), .D(
        n837), .Y(n817) );
  NOR2X1 U421 ( .A(n938), .B(n937), .Y(n941) );
  OAI31X1 U422 ( .A0(n938), .A1(n937), .A2(n2761), .B0(n936), .Y(n954) );
  OA21X1 U423 ( .A0(n921), .A1(n920), .B0(n919), .Y(n937) );
  NOR2X1 U424 ( .A(n503), .B(n502), .Y(n501) );
  CLKINVX1 U425 ( .A(n2188), .Y(n2209) );
  OA21X2 U426 ( .A0(n2556), .A1(n2557), .B0(n2555), .Y(n2567) );
  CLKINVX1 U427 ( .A(n2552), .Y(n2556) );
  NAND2X1 U428 ( .A(n2392), .B(n2404), .Y(n2400) );
  NAND2X1 U429 ( .A(n384), .B(n1556), .Y(n1786) );
  XOR2X1 U430 ( .A(\intadd_3/A[9] ), .B(n245), .Y(\intadd_3/SUM[9] ) );
  AND2X2 U431 ( .A(\intadd_3/B[8] ), .B(\intadd_3/n3 ), .Y(n245) );
  CLKINVX1 U432 ( .A(n310), .Y(n1917) );
  AOI2BB1X2 U433 ( .A0N(cr_read_cntr[6]), .A1N(n2703), .B0(n1025), .Y(n1030)
         );
  AOI32X1 U434 ( .A0(cr_read_cntr[6]), .A1(n1024), .A2(n2703), .B0(n301), .B1(
        n1023), .Y(n1026) );
  NAND2X1 U435 ( .A(cr_read_cntr[7]), .B(n225), .Y(n2703) );
  NOR2X1 U436 ( .A(n860), .B(n859), .Y(n853) );
  CLKINVX1 U437 ( .A(n850), .Y(n860) );
  OAI21X1 U438 ( .A0(n2289), .A1(n2280), .B0(n2257), .Y(n2258) );
  NAND2X1 U439 ( .A(n2254), .B(n2264), .Y(n2280) );
  NAND2X1 U440 ( .A(n2278), .B(n2294), .Y(n2267) );
  NOR2X1 U441 ( .A(n2255), .B(n2280), .Y(n2278) );
  OAI21X1 U442 ( .A0(n1440), .A1(n1433), .B0(n2423), .Y(n1434) );
  NAND2BX1 U443 ( .AN(n1440), .B(n1439), .Y(n1443) );
  NOR2X1 U444 ( .A(n1432), .B(n1431), .Y(n1440) );
  NAND2X1 U445 ( .A(next_state[1]), .B(n17), .Y(n1894) );
  NAND2X1 U446 ( .A(n316), .B(n232), .Y(n2102) );
  INVX4 U447 ( .A(n317), .Y(n316) );
  OAI31X1 U448 ( .A0(n2661), .A1(n138), .A2(n2660), .B0(n2659), .Y(n2666) );
  NAND2X1 U449 ( .A(n2651), .B(n2653), .Y(n2661) );
  CLKINVX1 U450 ( .A(n554), .Y(n540) );
  AOI211X1 U451 ( .A0(n1726), .A1(n1731), .B0(n1724), .C0(n1728), .Y(n1727) );
  NAND2X1 U452 ( .A(n1715), .B(n1714), .Y(n1731) );
  CLKINVX1 U453 ( .A(n1551), .Y(n1278) );
  NOR2X1 U454 ( .A(n2167), .B(n2166), .Y(n2168) );
  AND2X2 U455 ( .A(n2185), .B(n2181), .Y(n2166) );
  OAI21X1 U456 ( .A0(n1268), .A1(n1267), .B0(n1266), .Y(n1269) );
  NAND2X1 U457 ( .A(n232), .B(n1236), .Y(n1267) );
  NOR2X1 U458 ( .A(n1258), .B(n1267), .Y(n1257) );
  NOR2BX1 U459 ( .AN(n1262), .B(n1258), .Y(n1265) );
  OAI31X1 U460 ( .A0(n1226), .A1(n1258), .A2(n1225), .B0(n1231), .Y(n1261) );
  NAND2X1 U461 ( .A(n1270), .B(n1279), .Y(n1258) );
  NOR2X1 U462 ( .A(work_cntr[19]), .B(n2388), .Y(n2391) );
  CLKINVX1 U463 ( .A(n1812), .Y(n2774) );
  NAND2X1 U464 ( .A(n948), .B(n950), .Y(n956) );
  NAND2X1 U465 ( .A(n2243), .B(n2242), .Y(n2244) );
  AOI2BB2X2 U466 ( .B0(n2113), .B1(n2127), .A0N(n2113), .A1N(n2127), .Y(n2140)
         );
  NAND2X1 U467 ( .A(n2128), .B(n130), .Y(n2127) );
  NAND2X1 U468 ( .A(n1604), .B(n1798), .Y(n1610) );
  NOR2X1 U469 ( .A(n2232), .B(n2260), .Y(n2256) );
  NOR2X1 U470 ( .A(n1782), .B(n318), .Y(expand_sel[3]) );
  NAND2X1 U471 ( .A(n2008), .B(n2007), .Y(n2019) );
  AOI2BB2X2 U472 ( .B0(next_work_cntr[11]), .B1(n1998), .A0N(
        next_work_cntr[11]), .A1N(n1998), .Y(n2008) );
  NOR2X1 U473 ( .A(curr_time[1]), .B(n512), .Y(n510) );
  NOR2X1 U474 ( .A(n1866), .B(n1865), .Y(n1861) );
  NAND2X1 U475 ( .A(n1420), .B(n1421), .Y(n1415) );
  OA21X1 U476 ( .A0(n901), .A1(n900), .B0(n899), .Y(n911) );
  NAND2X1 U477 ( .A(n1402), .B(n1771), .Y(n2812) );
  OAI21X1 U478 ( .A0(n916), .A1(n915), .B0(n914), .Y(n918) );
  CLKINVX1 U479 ( .A(n2812), .Y(n2873) );
  NAND2BX1 U480 ( .AN(n912), .B(n911), .Y(n915) );
  NAND2X1 U481 ( .A(n921), .B(n1880), .Y(n922) );
  CLKINVX1 U482 ( .A(n2294), .Y(n2277) );
  NOR2X1 U483 ( .A(n2872), .B(n284), .Y(n2862) );
  CLKINVX1 U484 ( .A(n747), .Y(n1787) );
  NOR2BX1 U485 ( .AN(n2521), .B(n2119), .Y(n2114) );
  OAI22X1 U486 ( .A0(n1875), .A1(n1874), .B0(n1873), .B1(n1936), .Y(n1876) );
  NOR2X1 U487 ( .A(n1855), .B(n1932), .Y(n1875) );
  OAI2BB2X2 U488 ( .B0(n1187), .B1(n1186), .A0N(n1187), .A1N(n1186), .Y(n1235)
         );
  NAND2X1 U489 ( .A(n1185), .B(n1214), .Y(n1186) );
  OAI21X1 U490 ( .A0(n1495), .A1(n1490), .B0(n264), .Y(n1496) );
  NOR2BX1 U491 ( .AN(n1483), .B(n1482), .Y(n1490) );
  NOR2X1 U492 ( .A(work_cntr[19]), .B(n2386), .Y(n2514) );
  OAI21X1 U493 ( .A0(n2417), .A1(n251), .B0(n2416), .Y(n2431) );
  NOR2X1 U494 ( .A(work_cntr[10]), .B(n2433), .Y(n2417) );
  CLKINVX1 U495 ( .A(n2136), .Y(n2143) );
  NOR2X1 U496 ( .A(n2143), .B(n2138), .Y(n2193) );
  NOR2X1 U497 ( .A(n1653), .B(n1659), .Y(n1647) );
  CLKINVX1 U498 ( .A(n1665), .Y(n1659) );
  NAND3X1 U499 ( .A(n1832), .B(n1018), .C(n877), .Y(n1012) );
  OAI31X1 U500 ( .A0(n1993), .A1(n1990), .A2(n1984), .B0(n1983), .Y(n1987) );
  NOR2X1 U501 ( .A(n1980), .B(n1992), .Y(n1990) );
  NAND2X1 U502 ( .A(n1620), .B(write_cntr[7]), .Y(n1585) );
  CLKINVX1 U503 ( .A(n1583), .Y(n1620) );
  NOR2X1 U504 ( .A(n2315), .B(n2309), .Y(n2279) );
  NAND2X1 U505 ( .A(n1577), .B(n1620), .Y(n1582) );
  NAND3X1 U506 ( .A(n2343), .B(n2337), .C(n2355), .Y(n2347) );
  NOR2X1 U507 ( .A(n2320), .B(n2341), .Y(n2355) );
  NOR2BX1 U508 ( .AN(n824), .B(n1938), .Y(n825) );
  NOR2X2 U509 ( .A(n2766), .B(n2765), .Y(n2773) );
  OAI21X1 U510 ( .A0(n1586), .A1(n1585), .B0(n1584), .Y(n1587) );
  AOI21X1 U511 ( .A0(n1567), .A1(n1584), .B0(n1566), .Y(n1568) );
  NAND2X1 U512 ( .A(write_cntr[8]), .B(n1621), .Y(n1584) );
  NOR2X1 U513 ( .A(n1071), .B(n1051), .Y(n1049) );
  NAND2BX1 U514 ( .AN(n1605), .B(n1606), .Y(n1628) );
  NAND2X1 U515 ( .A(n287), .B(n1594), .Y(n1606) );
  CLKINVX1 U516 ( .A(n226), .Y(n2718) );
  NAND2BX1 U517 ( .AN(n1595), .B(n1619), .Y(n1599) );
  NOR2X1 U518 ( .A(n2216), .B(n2221), .Y(n2225) );
  NOR2X1 U519 ( .A(n1241), .B(n1201), .Y(n1219) );
  NOR2X1 U520 ( .A(n2122), .B(n2125), .Y(n2123) );
  NOR2X1 U521 ( .A(n2582), .B(n2115), .Y(n2122) );
  NOR2X1 U522 ( .A(n2227), .B(n2226), .Y(n2234) );
  NAND2X1 U523 ( .A(n2295), .B(n2294), .Y(n2318) );
  NOR2X1 U524 ( .A(n1605), .B(n1625), .Y(n1607) );
  NOR2X1 U525 ( .A(n1622), .B(n274), .Y(n1625) );
  NOR2X1 U526 ( .A(n1084), .B(n1082), .Y(n1121) );
  NAND2X1 U527 ( .A(global_cntr[7]), .B(n326), .Y(n327) );
  NAND2X1 U528 ( .A(n2039), .B(n2040), .Y(n1957) );
  NAND2X1 U529 ( .A(n316), .B(n2620), .Y(n2039) );
  NOR2X1 U530 ( .A(n1121), .B(n1120), .Y(n1123) );
  NAND2BX1 U531 ( .AN(n2333), .B(n2332), .Y(n2364) );
  NOR2X1 U532 ( .A(n235), .B(n2829), .Y(n1814) );
  NAND2X1 U533 ( .A(curr_time[23]), .B(n972), .Y(n431) );
  NAND2X1 U534 ( .A(global_cntr[9]), .B(n328), .Y(n332) );
  NOR2BX1 U535 ( .AN(n1012), .B(n1933), .Y(n1013) );
  CLKINVX1 U536 ( .A(n306), .Y(n2681) );
  NOR2X1 U537 ( .A(n2131), .B(n2130), .Y(n2132) );
  NOR2X1 U538 ( .A(n2277), .B(n2298), .Y(n2266) );
  NOR2X1 U539 ( .A(n283), .B(n2776), .Y(n2779) );
  NOR2X1 U540 ( .A(n2075), .B(n2078), .Y(n2090) );
  NOR2X1 U541 ( .A(n2068), .B(n2067), .Y(n2075) );
  NOR2X1 U542 ( .A(n1099), .B(n1126), .Y(n1130) );
  NOR2BX1 U543 ( .AN(n1104), .B(n1125), .Y(n1099) );
  NOR2BX1 U544 ( .AN(n1833), .B(n1925), .Y(n1835) );
  NOR2X1 U545 ( .A(n1039), .B(n1412), .Y(n1059) );
  AOI21X1 U546 ( .A0(n1161), .A1(n1159), .B0(n1167), .Y(n1165) );
  NOR2X1 U547 ( .A(n1168), .B(n1197), .Y(n1161) );
  NOR2BX1 U548 ( .AN(n1205), .B(n1194), .Y(n1193) );
  NOR2BX1 U549 ( .AN(n1204), .B(n1195), .Y(n1194) );
  OAI21X1 U550 ( .A0(n1106), .A1(n1129), .B0(n1105), .Y(n1107) );
  NAND2X1 U551 ( .A(n1126), .B(n1099), .Y(n1129) );
  NOR2BX1 U552 ( .AN(n1430), .B(n1428), .Y(n1433) );
  NOR2X1 U553 ( .A(n1427), .B(n1419), .Y(n1428) );
  NAND2BX1 U554 ( .AN(n1229), .B(n1227), .Y(n1212) );
  AOI21X1 U555 ( .A0(n1195), .A1(n1205), .B0(n1194), .Y(n1229) );
  NOR2X1 U556 ( .A(n1933), .B(n1932), .Y(n1943) );
  NOR2BX1 U557 ( .AN(n1524), .B(n1519), .Y(n1527) );
  NOR2X1 U558 ( .A(cr_read_cntr[5]), .B(n1026), .Y(n1028) );
  NOR2X1 U559 ( .A(n1938), .B(n1937), .Y(n2705) );
  NOR3X1 U560 ( .A(work_cntr[4]), .B(n2074), .C(n317), .Y(n2078) );
  NOR2X1 U561 ( .A(n2066), .B(n2067), .Y(n2074) );
  OAI21X1 U562 ( .A0(n2817), .A1(n2853), .B0(n2851), .Y(n2856) );
  NOR2BX1 U563 ( .AN(n1662), .B(n1676), .Y(n1678) );
  NAND2X1 U564 ( .A(write_addr[15]), .B(write_addr[14]), .Y(n1812) );
  NOR2BX1 U565 ( .AN(n1670), .B(n1669), .Y(n1673) );
  OAI21X1 U566 ( .A0(n1678), .A1(n1668), .B0(n1667), .Y(n1670) );
  NAND2X1 U567 ( .A(n1832), .B(n1830), .Y(n1833) );
  NOR2BX1 U568 ( .AN(n1850), .B(n1848), .Y(n1830) );
  NAND2BX1 U569 ( .AN(n1543), .B(n232), .Y(n1538) );
  OAI21X1 U570 ( .A0(n1534), .A1(n263), .B0(n1533), .Y(n1543) );
  NAND2BX1 U571 ( .AN(n1067), .B(n2423), .Y(n1072) );
  NOR2X1 U572 ( .A(n1996), .B(n1997), .Y(n2003) );
  AOI31X1 U573 ( .A0(n2004), .A1(n1995), .A2(n1994), .B0(n1993), .Y(n1996) );
  NAND2X1 U574 ( .A(n2079), .B(n2068), .Y(n2071) );
  OAI2BB2X1 U575 ( .B0(n1347), .B1(n1346), .A0N(n1347), .A1N(n1345), .Y(n1351)
         );
  OAI21X1 U576 ( .A0(n1343), .A1(n1342), .B0(n1341), .Y(n1347) );
  NOR3X1 U577 ( .A(n2820), .B(n296), .C(n224), .Y(n2822) );
  OAI21X1 U578 ( .A0(n1101), .A1(n1109), .B0(n1100), .Y(n1102) );
  NAND2X1 U579 ( .A(n1889), .B(n1886), .Y(n1926) );
  OAI21X1 U580 ( .A0(n1872), .A1(n1871), .B0(n1870), .Y(n1886) );
  NOR2X1 U581 ( .A(n1516), .B(n1515), .Y(n1519) );
  OAI21X1 U582 ( .A0(n1509), .A1(n1513), .B0(n1508), .Y(n1515) );
  NOR2X1 U583 ( .A(n1937), .B(n1922), .Y(n1935) );
  OAI21X1 U584 ( .A0(n1921), .A1(n1920), .B0(n1919), .Y(n1922) );
  NOR3X1 U585 ( .A(n2791), .B(n2790), .C(n2789), .Y(n2792) );
  NOR3X1 U586 ( .A(n2789), .B(n1639), .C(N2294), .Y(en_fb_addr) );
  CLKINVX1 U587 ( .A(n769), .Y(n2789) );
  OAI21X1 U588 ( .A0(n1536), .A1(n1535), .B0(n232), .Y(n1542) );
  AOI22X1 U589 ( .A0(n1390), .A1(n1389), .B0(n1388), .B1(n1387), .Y(n1394) );
  OAI21X1 U590 ( .A0(n1386), .A1(n1385), .B0(n1384), .Y(n1390) );
  NAND2X1 U591 ( .A(n2326), .B(n2344), .Y(n2327) );
  OAI21X1 U592 ( .A0(n2325), .A1(n2324), .B0(n2323), .Y(n2344) );
  NOR2X1 U593 ( .A(n1661), .B(n1660), .Y(n1674) );
  OAI21X1 U594 ( .A0(n1654), .A1(n1653), .B0(n1652), .Y(n1661) );
  OAI21X1 U595 ( .A0(n2349), .A1(n2348), .B0(n2358), .Y(n2350) );
  OAI21X1 U596 ( .A0(n2347), .A1(n2346), .B0(n2345), .Y(n2358) );
  OAI211X1 U597 ( .A0(n2506), .A1(n2507), .B0(n2505), .C0(n2504), .Y(n2511) );
  NOR2X1 U598 ( .A(n1480), .B(n1479), .Y(n1482) );
  OAI21X1 U599 ( .A0(n140), .A1(n1477), .B0(n1472), .Y(n1480) );
  OAI211X1 U600 ( .A0(n545), .A1(n553), .B0(n544), .C0(n543), .Y(\C1/Z_0 ) );
  NOR2X1 U601 ( .A(n285), .B(n2802), .Y(n738) );
  NOR2X1 U602 ( .A(n2807), .B(n285), .Y(n2842) );
  OAI2BB2X1 U603 ( .B0(next_work_cntr[17]), .B1(n2132), .A0N(
        next_work_cntr[17]), .A1N(n2132), .Y(n2162) );
  AOI211X4 U604 ( .A0(n2684), .A1(n310), .B0(n2683), .C0(n744), .Y(n2690) );
  NAND3X1 U605 ( .A(n805), .B(n808), .C(n806), .Y(n2684) );
  OAI21X1 U606 ( .A0(n1522), .A1(n1523), .B0(n1521), .Y(n1525) );
  OAI21X1 U607 ( .A0(n1727), .A1(n1722), .B0(n1721), .Y(n1725) );
  NOR2X1 U608 ( .A(n1036), .B(work_cntr[10]), .Y(n1043) );
  OAI21X1 U609 ( .A0(n1059), .A1(n1058), .B0(n1057), .Y(n1087) );
  OAI21X2 U610 ( .A0(n1283), .A1(n1401), .B0(work_cntr[19]), .Y(n1036) );
  NOR3X1 U611 ( .A(next_work_cntr[4]), .B(n2309), .C(n2263), .Y(n2254) );
  CLKINVX1 U612 ( .A(n2225), .Y(n2263) );
  AOI2BB2X2 U613 ( .B0(n166), .B1(n2230), .A0N(n166), .A1N(n2230), .Y(n2238)
         );
  OAI21X1 U614 ( .A0(n2229), .A1(n2234), .B0(n2228), .Y(n2230) );
  AOI2BB2X2 U615 ( .B0(n2263), .B1(n2262), .A0N(n2263), .A1N(n2262), .Y(n2315)
         );
  OAI21X1 U616 ( .A0(n2261), .A1(n2283), .B0(n2260), .Y(n2262) );
  OAI21X1 U617 ( .A0(n1130), .A1(n1155), .B0(n1129), .Y(n1131) );
  OAI21X1 U618 ( .A0(n2810), .A1(n2803), .B0(n2800), .Y(n2841) );
  AOI21X1 U619 ( .A0(n2304), .A1(n2303), .B0(n2302), .Y(n2324) );
  OAI2BB2X1 U620 ( .B0(n2269), .B1(n2268), .A0N(n2269), .A1N(n2268), .Y(n2304)
         );
  OAI21X1 U621 ( .A0(n1425), .A1(n1429), .B0(n1424), .Y(n1431) );
  OAI21X1 U622 ( .A0(n1428), .A1(n1423), .B0(n216), .Y(n1429) );
  CLKINVX1 U623 ( .A(n1098), .Y(n1126) );
  NOR3X2 U624 ( .A(n1098), .B(n1132), .C(n1086), .Y(n1096) );
  AOI22X1 U625 ( .A0(n1070), .A1(work_cntr[13]), .B0(n1069), .B1(n1068), .Y(
        n1098) );
  OAI2BB2X1 U626 ( .B0(n1241), .B1(n1240), .A0N(n1241), .A1N(n1240), .Y(n1274)
         );
  NOR2X1 U627 ( .A(n2054), .B(n2055), .Y(n2059) );
  OAI21X1 U628 ( .A0(n2052), .A1(n2051), .B0(n2050), .Y(n2055) );
  NOR2X1 U629 ( .A(n1768), .B(n232), .Y(n1776) );
  NAND3X1 U630 ( .A(write_addr[2]), .B(write_addr[1]), .C(write_addr[3]), .Y(
        n2837) );
  OAI21X1 U631 ( .A0(n1936), .A1(n1873), .B0(n1860), .Y(n1879) );
  NAND2X1 U632 ( .A(n316), .B(n830), .Y(n838) );
  NAND3X1 U633 ( .A(write_cntr[7]), .B(write_cntr[6]), .C(n837), .Y(n830) );
  NAND4X1 U634 ( .A(n228), .B(n251), .C(n217), .D(n2423), .Y(n1642) );
  NAND2X1 U635 ( .A(n1061), .B(n1074), .Y(n1105) );
  NOR2X1 U636 ( .A(work_cntr[13]), .B(n1066), .Y(n1074) );
  OAI22X1 U637 ( .A0(n2517), .A1(n2521), .B0(n2516), .B1(n259), .Y(n2523) );
  NOR2X1 U638 ( .A(n2411), .B(n2413), .Y(n2422) );
  OAI22X1 U639 ( .A0(n2421), .A1(n2410), .B0(n2409), .B1(n2408), .Y(n2413) );
  NOR2X1 U640 ( .A(n1039), .B(n1036), .Y(n1063) );
  OAI21X1 U641 ( .A0(n1216), .A1(n1266), .B0(n1215), .Y(n1217) );
  NOR2BX1 U642 ( .AN(n1193), .B(n273), .Y(n1216) );
  NOR3X1 U643 ( .A(write_addr[17]), .B(write_addr[18]), .C(n2797), .Y(n2806)
         );
  CLKINVX1 U644 ( .A(n1800), .Y(n743) );
  OR2X2 U645 ( .A(n1623), .B(n1638), .Y(n1800) );
  CLKINVX1 U646 ( .A(n2450), .Y(n2444) );
  OAI21X1 U647 ( .A0(n881), .A1(n880), .B0(n879), .Y(n887) );
  NOR3X1 U648 ( .A(n131), .B(n1879), .C(n1880), .Y(n1868) );
  NOR2X1 U649 ( .A(n275), .B(n833), .Y(n836) );
  NOR2X1 U650 ( .A(n1807), .B(n827), .Y(n828) );
  OAI22X1 U651 ( .A0(n1011), .A1(n1010), .B0(n1019), .B1(n1009), .Y(n1838) );
  AOI211X4 U652 ( .A0(n1278), .A1(n1277), .B0(n1276), .C0(n1275), .Y(n1557) );
  NAND2BX1 U653 ( .AN(n2302), .B(n2303), .Y(n2290) );
  NOR3X1 U654 ( .A(next_work_cntr[16]), .B(next_work_cntr[17]), .C(n2124), .Y(
        n2118) );
  AOI211X1 U655 ( .A0(n263), .A1(n1756), .B0(n1762), .C0(n1755), .Y(n1767) );
  OAI21X1 U656 ( .A0(next_en_si), .A1(n317), .B0(n2771), .Y(n2683) );
  OAI22X2 U657 ( .A0(n2709), .A1(n2680), .B0(n2679), .B1(n2783), .Y(next_en_si) );
  NOR2X1 U658 ( .A(n1761), .B(n1760), .Y(n1777) );
  NOR3X1 U659 ( .A(n273), .B(n1755), .C(n1759), .Y(n1761) );
  OAI2BB2X1 U660 ( .B0(n2343), .B1(n2342), .A0N(n2343), .A1N(n2342), .Y(n2362)
         );
  OAI31X1 U661 ( .A0(n2341), .A1(n2340), .A2(n2339), .B0(n2338), .Y(n2342) );
  OAI21X1 U662 ( .A0(n1761), .A1(n1754), .B0(N1827), .Y(n1756) );
  NOR2X1 U663 ( .A(N1827), .B(n1754), .Y(n1762) );
  OAI31X1 U664 ( .A0(n1753), .A1(n1752), .A2(n1751), .B0(n1750), .Y(n1754) );
  OAI21X1 U665 ( .A0(n1090), .A1(n1089), .B0(n1088), .Y(n1095) );
  NAND2X1 U666 ( .A(n1088), .B(n1087), .Y(n1085) );
  OAI21X1 U667 ( .A0(n1147), .A1(n1146), .B0(n1145), .Y(n1166) );
  OAI31X1 U668 ( .A0(n1134), .A1(n1133), .A2(n1138), .B0(n1147), .Y(n1145) );
  OAI31X1 U669 ( .A0(n2098), .A1(n2097), .A2(n2096), .B0(n2095), .Y(n2103) );
  OAI21X1 U670 ( .A0(n2038), .A1(n2046), .B0(n2037), .Y(n2041) );
  AOI221X1 U671 ( .A0(n2044), .A1(n2036), .B0(n2057), .B1(n2036), .C0(n2043), 
        .Y(n2046) );
  NOR2X1 U672 ( .A(N196), .B(n1552), .Y(n1262) );
  NOR2X1 U673 ( .A(n1552), .B(n2863), .Y(n1556) );
  AOI2BB2X2 U674 ( .B0(N1825), .B1(n1236), .A0N(N1825), .A1N(n1236), .Y(n1552)
         );
  OAI21X1 U675 ( .A0(n1197), .A1(n1210), .B0(n1196), .Y(n1200) );
  OAI21X1 U676 ( .A0(n2421), .A1(n2420), .B0(n2419), .Y(n2426) );
  NOR2X1 U677 ( .A(n2333), .B(n2365), .Y(n2354) );
  XOR2X1 U678 ( .A(n2311), .B(n2315), .Y(n2365) );
  NOR2X2 U679 ( .A(n232), .B(n284), .Y(n1789) );
  OAI21X1 U680 ( .A0(N1826), .A1(n1789), .B0(n2668), .Y(n1952) );
  XNOR2X1 U681 ( .A(read_cntr[0]), .B(read_cntr[1]), .Y(n2811) );
  NOR2BX1 U682 ( .AN(n2815), .B(n1789), .Y(n2859) );
  AOI2BB2X2 U683 ( .B0(n1018), .B1(n1017), .A0N(n1018), .A1N(n1017), .Y(n1834)
         );
  OAI21X1 U684 ( .A0(cr_read_cntr[7]), .A1(n2699), .B0(n2698), .Y(n2701) );
  AOI221X1 U685 ( .A0(n2696), .A1(n2695), .B0(n301), .B1(n2695), .C0(n2694), 
        .Y(n2698) );
  NOR3X1 U686 ( .A(n1988), .B(n169), .C(n1992), .Y(n1993) );
  AOI2BB2X2 U687 ( .B0(next_work_cntr[13]), .B1(n1985), .A0N(
        next_work_cntr[13]), .A1N(n1985), .Y(n1988) );
  AOI2BB2X2 U688 ( .B0(n310), .B1(\intadd_3/SUM[9] ), .A0N(n2764), .A1N(n2783), 
        .Y(n632) );
  NOR3BX1 U689 ( .AN(n1598), .B(n1595), .C(n1600), .Y(n1602) );
  AOI2BB2X2 U690 ( .B0(n310), .B1(\intadd_3/SUM[3] ), .A0N(n2839), .A1N(n776), 
        .Y(n2845) );
  AOI2BB2X2 U691 ( .B0(n1588), .B1(n1587), .A0N(n1588), .A1N(n1587), .Y(n1600)
         );
  AOI2BB2X2 U692 ( .B0(n136), .B1(n2018), .A0N(n136), .A1N(n2018), .Y(n2028)
         );
  OAI31X1 U693 ( .A0(n1704), .A1(n1703), .A2(n1702), .B0(n1701), .Y(n1708) );
  AOI2BB2X2 U694 ( .B0(n1683), .B1(n1685), .A0N(n1683), .A1N(n1685), .Y(n1702)
         );
  NOR4X1 U695 ( .A(global_cntr[7]), .B(global_cntr[8]), .C(global_cntr[15]), 
        .D(n777), .Y(n1553) );
  NOR4X1 U696 ( .A(n760), .B(n759), .C(n761), .D(n762), .Y(n795) );
  AOI2BB2X2 U697 ( .B0(work_cntr[19]), .B1(n2516), .A0N(work_cntr[19]), .A1N(
        n2516), .Y(n2522) );
  NOR2X2 U698 ( .A(n250), .B(n325), .Y(n758) );
  NAND2X1 U699 ( .A(n458), .B(n457), .Y(n513) );
  NOR2X1 U700 ( .A(n433), .B(n432), .Y(n457) );
  NOR2X1 U701 ( .A(next_work_cntr[8]), .B(n2143), .Y(n2185) );
  OAI2BB2X1 U702 ( .B0(n2129), .B1(n2159), .A0N(n2129), .A1N(
        next_work_cntr[15]), .Y(n2189) );
  NAND2X1 U703 ( .A(n2129), .B(n2128), .Y(n2139) );
  NOR2X1 U704 ( .A(n2157), .B(n2152), .Y(n2129) );
  NOR2BX1 U705 ( .AN(n2079), .B(n2077), .Y(n2083) );
  NOR2X1 U706 ( .A(N1827), .B(n317), .Y(n2077) );
  NOR2BX1 U707 ( .AN(n2205), .B(n2204), .Y(n2241) );
  NOR2BX1 U708 ( .AN(n2218), .B(n2220), .Y(n2204) );
  NOR2X1 U709 ( .A(n2315), .B(n2314), .Y(n2336) );
  OAI21X1 U710 ( .A0(n2831), .A1(n2853), .B0(n2851), .Y(n2832) );
  NOR2X1 U711 ( .A(n2829), .B(n281), .Y(n2831) );
  OAI22X1 U712 ( .A0(write_cntr[13]), .A1(n814), .B0(n279), .B1(n813), .Y(n841) );
  NOR2BX1 U713 ( .AN(n2493), .B(n2491), .Y(n2500) );
  NOR2X1 U714 ( .A(n265), .B(n815), .Y(n814) );
  OAI2BB2X1 U715 ( .B0(n1335), .B1(n1336), .A0N(n1335), .A1N(n1334), .Y(n1344)
         );
  NAND2X1 U716 ( .A(n2836), .B(write_addr[5]), .Y(n1818) );
  NOR2X1 U717 ( .A(n2837), .B(n741), .Y(n2836) );
  OAI21X1 U718 ( .A0(n1418), .A1(n1417), .B0(n1416), .Y(n1427) );
  NOR2X1 U719 ( .A(n2003), .B(n2010), .Y(n2012) );
  OAI2BB2X1 U720 ( .B0(n1410), .B1(n257), .A0N(n1410), .A1N(n257), .Y(n1418)
         );
  AOI2BB2X2 U721 ( .B0(n310), .B1(\intadd_3/SUM[2] ), .A0N(n776), .A1N(n2838), 
        .Y(n675) );
  OAI21X1 U722 ( .A0(n468), .A1(n467), .B0(n520), .Y(n541) );
  OAI21X1 U723 ( .A0(write_addr[5]), .A1(n2836), .B0(n1818), .Y(n2838) );
  OAI2BB2X1 U724 ( .B0(n2426), .B1(n2425), .A0N(n2426), .A1N(n2424), .Y(n2436)
         );
  OAI21X1 U725 ( .A0(n2436), .A1(n2435), .B0(n2434), .Y(n2440) );
  NOR2X1 U726 ( .A(n2689), .B(n302), .Y(n2692) );
  NAND3BX2 U727 ( .AN(n1008), .B(work_cntr[5]), .C(work_cntr[4]), .Y(n1948) );
  OAI211X1 U728 ( .A0(n1333), .A1(n1332), .B0(n1331), .C0(n1330), .Y(n1343) );
  CLKINVX1 U729 ( .A(n722), .Y(n703) );
  OAI211X1 U730 ( .A0(n2771), .A1(n288), .B0(n1904), .C0(n358), .Y(n722) );
  OAI21X1 U731 ( .A0(n228), .A1(n1463), .B0(n1462), .Y(n1467) );
  OAI21X1 U732 ( .A0(n2526), .A1(n2525), .B0(n2530), .Y(n2534) );
  AOI31X1 U733 ( .A0(n2709), .A1(n2708), .A2(n2707), .B0(n2706), .Y(n2846) );
  OAI21X1 U734 ( .A0(n273), .A1(n1524), .B0(n1523), .Y(n1530) );
  OAI21X1 U735 ( .A0(n1519), .A1(n1518), .B0(n273), .Y(n1523) );
  OAI21X1 U736 ( .A0(n1151), .A1(n1117), .B0(n1116), .Y(n1118) );
  NOR2BX1 U737 ( .AN(n172), .B(n1114), .Y(n1151) );
  OAI2BB2X2 U738 ( .B0(next_work_cntr[18]), .B1(n1960), .A0N(
        next_work_cntr[18]), .A1N(n1960), .Y(n1974) );
  NOR2BX1 U739 ( .AN(n1959), .B(next_work_cntr[17]), .Y(n1960) );
  AOI2BB2X2 U740 ( .B0(n1733), .B1(n212), .A0N(n1733), .A1N(n212), .Y(n1745)
         );
  NAND2X1 U741 ( .A(n1733), .B(n212), .Y(n1737) );
  NOR2X1 U742 ( .A(n885), .B(n886), .Y(n881) );
  OAI21X1 U743 ( .A0(n869), .A1(n868), .B0(n867), .Y(n885) );
  OAI21X1 U744 ( .A0(n2220), .A1(n2219), .B0(n2218), .Y(n2250) );
  AOI2BB1X2 U745 ( .A0N(n1672), .A1N(n2423), .B0(n1671), .Y(n1685) );
  NOR2X1 U746 ( .A(n1709), .B(n1642), .Y(n1671) );
  NOR2BX1 U747 ( .AN(n2061), .B(n2060), .Y(n2070) );
  OAI2BB2X1 U748 ( .B0(n2060), .B1(n2061), .A0N(n2060), .A1N(n2061), .Y(n2079)
         );
  OAI2BB2X1 U749 ( .B0(n1575), .B1(n1576), .A0N(n1575), .A1N(n1580), .Y(n1601)
         );
  OAI22X1 U750 ( .A0(n1565), .A1(n1564), .B0(n1563), .B1(n1572), .Y(n1575) );
  NOR2X1 U751 ( .A(work_cntr[9]), .B(n1045), .Y(n1044) );
  OAI21X1 U752 ( .A0(n1358), .A1(n1357), .B0(n1356), .Y(n1361) );
  OAI22X1 U753 ( .A0(n1339), .A1(n261), .B0(n1354), .B1(n1709), .Y(n1357) );
  NOR2X1 U754 ( .A(n1709), .B(n1283), .Y(n1644) );
  NOR2X1 U755 ( .A(n1367), .B(n1370), .Y(n1379) );
  CLKINVX1 U756 ( .A(n1367), .Y(n1375) );
  OAI22X1 U757 ( .A0(n1354), .A1(n1353), .B0(n1281), .B1(n264), .Y(n1367) );
  NOR3X2 U758 ( .A(n1124), .B(n1122), .C(n1119), .Y(n1104) );
  AOI2BB2X2 U759 ( .B0(n1084), .B1(n1083), .A0N(n1084), .A1N(n1083), .Y(n1119)
         );
  NAND2X1 U760 ( .A(n1002), .B(work_cntr[11]), .Y(n1001) );
  NOR2X1 U761 ( .A(n1003), .B(n228), .Y(n1002) );
  OAI31X1 U762 ( .A0(n892), .A1(n891), .A2(n890), .B0(n889), .Y(n905) );
  NAND2X1 U763 ( .A(n891), .B(n882), .Y(n896) );
  OAI22X1 U764 ( .A0(n877), .A1(n876), .B0(n875), .B1(n874), .Y(n891) );
  OAI22X1 U765 ( .A0(n1581), .A1(n1580), .B0(n1579), .B1(n1578), .Y(n1603) );
  OAI2BB2X2 U766 ( .B0(n894), .B1(n893), .A0N(n894), .A1N(n893), .Y(n907) );
  NOR2X1 U767 ( .A(n1873), .B(n913), .Y(n912) );
  OAI22X1 U768 ( .A0(n1857), .A1(n2742), .B0(n1846), .B1(n2737), .Y(n913) );
  OAI22X1 U769 ( .A0(n233), .A1(n2721), .B0(n2722), .B1(n2723), .Y(n2726) );
  AOI22X1 U770 ( .A0(n944), .A1(n943), .B0(n949), .B1(n953), .Y(n959) );
  OAI21X1 U771 ( .A0(n941), .A1(n940), .B0(n939), .Y(n949) );
  INVXL U772 ( .A(n1320), .Y(n156) );
  CLKINVX1 U773 ( .A(n156), .Y(n157) );
  OAI22X1 U774 ( .A0(n1864), .A1(n1863), .B0(n1869), .B1(n1862), .Y(n1887) );
  OAI21X1 U775 ( .A0(n1854), .A1(n1853), .B0(n1852), .Y(n1869) );
  OAI22X1 U776 ( .A0(n1828), .A1(n1827), .B0(n1836), .B1(n1826), .Y(n1853) );
  OAI21X1 U777 ( .A0(n1022), .A1(n1021), .B0(n1020), .Y(n1836) );
  OAI22X1 U778 ( .A0(n1842), .A1(n1841), .B0(n1851), .B1(n1840), .Y(n1871) );
  OAI21X1 U779 ( .A0(n1839), .A1(n1838), .B0(n1837), .Y(n1851) );
  OAI2BB2X1 U780 ( .B0(n2259), .B1(n2258), .A0N(n2259), .A1N(n2258), .Y(n2288)
         );
  AOI2BB2X2 U781 ( .B0(n2203), .B1(n2202), .A0N(n2203), .A1N(n2202), .Y(n2259)
         );
  OAI22X2 U782 ( .A0(N1825), .A1(N196), .B0(n232), .B1(n284), .Y(n2664) );
  AOI2BB2X2 U783 ( .B0(next_work_cntr[17]), .B1(n1959), .A0N(
        next_work_cntr[17]), .A1N(n1959), .Y(n1970) );
  AOI2BB2X2 U784 ( .B0(n2115), .B1(next_work_cntr[10]), .A0N(n2115), .A1N(
        n2582), .Y(n2169) );
  CLKINVX1 U785 ( .A(n2778), .Y(n158) );
  CLKINVX1 U786 ( .A(n158), .Y(n159) );
  OAI21X1 U787 ( .A0(n897), .A1(n896), .B0(n895), .Y(n898) );
  AOI2BB2X2 U788 ( .B0(work_cntr[15]), .B1(n1298), .A0N(work_cntr[15]), .A1N(
        n1298), .Y(n1308) );
  NOR2X1 U789 ( .A(work_cntr[14]), .B(n1312), .Y(n1298) );
  NOR3X2 U790 ( .A(N1826), .B(n317), .C(n2084), .Y(n2100) );
  CLKINVX1 U791 ( .A(n926), .Y(n160) );
  CLKINVX1 U792 ( .A(n160), .Y(n161) );
  OAI31X1 U793 ( .A0(n2158), .A1(n2157), .A2(n2176), .B0(n2156), .Y(n2188) );
  AND2X2 U794 ( .A(n2155), .B(n2190), .Y(n2176) );
  AOI2BB2X2 U795 ( .B0(n1175), .B1(n1176), .A0N(n1175), .A1N(n1176), .Y(n1221)
         );
  OAI31X4 U796 ( .A0(n1151), .A1(n1154), .A2(n1153), .B0(n1150), .Y(n1175) );
  OAI2BB2X1 U797 ( .B0(n270), .B1(n1749), .A0N(n270), .A1N(n1749), .Y(n1765)
         );
  INVXL U798 ( .A(n934), .Y(n162) );
  CLKINVX1 U799 ( .A(n162), .Y(n163) );
  NOR2BX1 U800 ( .AN(n2312), .B(n2331), .Y(n2308) );
  AOI2BB2X2 U801 ( .B0(next_work_cntr[3]), .B1(n2290), .A0N(next_work_cntr[3]), 
        .A1N(n2290), .Y(n2331) );
  OAI21X1 U802 ( .A0(n2545), .A1(n2544), .B0(n2547), .Y(n2551) );
  NAND3X1 U803 ( .A(n2581), .B(n2545), .C(n2556), .Y(n2112) );
  OAI21X2 U804 ( .A0(n998), .A1(work_cntr[14]), .B0(n997), .Y(n2545) );
  AOI2BB1X2 U805 ( .A0N(n970), .A1N(n963), .B0(n967), .Y(n2710) );
  OAI31X4 U806 ( .A0(n957), .A1(n2717), .A2(n956), .B0(n955), .Y(n967) );
  CLKINVX1 U807 ( .A(n737), .Y(n719) );
  OAI21X2 U808 ( .A0(n1311), .A1(n217), .B0(n1310), .Y(n1329) );
  CLKINVX1 U809 ( .A(n2482), .Y(n164) );
  NOR2X1 U810 ( .A(n264), .B(n1127), .Y(n1140) );
  NAND2X1 U811 ( .A(n264), .B(n1127), .Y(n1139) );
  NAND2X1 U812 ( .A(n1113), .B(n1127), .Y(n1114) );
  NAND2BX1 U813 ( .AN(n1136), .B(n1135), .Y(n1127) );
  OAI2BB2X1 U814 ( .B0(n907), .B1(n906), .A0N(n907), .A1N(n906), .Y(n916) );
  OAI22X1 U815 ( .A0(n1063), .A1(n257), .B0(n1283), .B1(n2515), .Y(n1051) );
  NAND2X1 U816 ( .A(work_cntr[19]), .B(n1401), .Y(n2515) );
  NAND2BX1 U817 ( .AN(n1734), .B(n1729), .Y(n1738) );
  NOR2X1 U818 ( .A(n1174), .B(n1191), .Y(n1160) );
  OAI2BB2X2 U819 ( .B0(n1174), .B1(n1173), .A0N(n1174), .A1N(n1173), .Y(n1187)
         );
  NAND2BX1 U820 ( .AN(n1140), .B(n1139), .Y(n1174) );
  NAND2BX1 U821 ( .AN(n1186), .B(n1187), .Y(n1232) );
  OAI2BB2X1 U822 ( .B0(curr_time[4]), .B1(\s_1[3] ), .A0N(curr_time[4]), .A1N(
        \s_1[3] ), .Y(n991) );
  NAND2X1 U823 ( .A(n349), .B(n353), .Y(\s_1[3] ) );
  NOR2X1 U824 ( .A(n424), .B(n547), .Y(n550) );
  OAI21X1 U825 ( .A0(n1671), .A1(n216), .B0(n1655), .Y(n1669) );
  CLKINVX1 U826 ( .A(n1655), .Y(n2382) );
  OAI22X1 U827 ( .A0(work_cntr[15]), .A1(n1655), .B0(n227), .B1(n2382), .Y(
        n1660) );
  NAND2X1 U828 ( .A(n1671), .B(n216), .Y(n1655) );
  NOR3X1 U829 ( .A(work_cntr[8]), .B(n1079), .C(n1103), .Y(n1060) );
  NOR2X1 U830 ( .A(n1103), .B(n1112), .Y(n1097) );
  NAND2X1 U831 ( .A(n1076), .B(n1075), .Y(n1103) );
  NOR2BX2 U832 ( .AN(n2306), .B(n2275), .Y(n2295) );
  NOR2X2 U833 ( .A(n410), .B(n548), .Y(n551) );
  NOR3X1 U834 ( .A(next_work_cntr[6]), .B(n2227), .C(n2217), .Y(n2205) );
  NOR2X1 U835 ( .A(next_work_cntr[6]), .B(n2204), .Y(n2216) );
  CLKINVX1 U836 ( .A(n2039), .Y(next_work_cntr[6]) );
  NOR2X1 U837 ( .A(n1621), .B(write_cntr[8]), .Y(n1586) );
  NAND2X1 U838 ( .A(n1562), .B(n1621), .Y(n1569) );
  NOR4X1 U839 ( .A(n1621), .B(n1620), .C(n1619), .D(n277), .Y(n1799) );
  OAI21X1 U840 ( .A0(n1081), .A1(n2381), .B0(n1080), .Y(n1122) );
  NOR2X1 U841 ( .A(n2381), .B(n1079), .Y(n1040) );
  AOI221X1 U842 ( .A0(n2381), .A1(work_cntr[13]), .B0(n1034), .B1(
        work_cntr[13]), .C0(n1035), .Y(n1068) );
  NAND2X1 U843 ( .A(n251), .B(n217), .Y(n2381) );
  OAI21X2 U844 ( .A0(work_cntr[5]), .A1(n1007), .B0(n1948), .Y(n2634) );
  NOR2X1 U845 ( .A(n270), .B(n1008), .Y(n1007) );
  OAI21X2 U846 ( .A0(n2447), .A1(n261), .B0(n2433), .Y(n2453) );
  NAND2X1 U847 ( .A(n2447), .B(n261), .Y(n2433) );
  NOR2X1 U848 ( .A(n2477), .B(n2380), .Y(n2447) );
  NAND2X1 U849 ( .A(n1708), .B(n1716), .Y(n1719) );
  AOI21X2 U850 ( .A0(n999), .A1(n2423), .B0(n998), .Y(n2552) );
  NOR2X1 U851 ( .A(n999), .B(n2423), .Y(n998) );
  OAI21X1 U852 ( .A0(n847), .A1(n846), .B0(n845), .Y(n859) );
  CLKINVX1 U853 ( .A(n840), .Y(n847) );
  OAI21X2 U854 ( .A0(n1387), .A1(n1382), .B0(n1389), .Y(n1393) );
  OAI21X1 U855 ( .A0(n1381), .A1(n1382), .B0(n1387), .Y(n1389) );
  OAI22X1 U856 ( .A0(n1386), .A1(n1380), .B0(n1379), .B1(n1378), .Y(n1382) );
  NAND2X1 U857 ( .A(n284), .B(n316), .Y(n2351) );
  OAI2BB2X1 U858 ( .B0(n2236), .B1(n2235), .A0N(n2236), .A1N(n2235), .Y(n2294)
         );
  NAND2X1 U859 ( .A(n2187), .B(n2228), .Y(n2236) );
  OAI21X1 U860 ( .A0(n2237), .A1(n2195), .B0(n2219), .Y(n2218) );
  NOR2BX1 U861 ( .AN(n2241), .B(n2237), .Y(n2210) );
  CLKINVX1 U862 ( .A(n2237), .Y(n2243) );
  OAI31X4 U863 ( .A0(n2173), .A1(n2172), .A2(n2175), .B0(n2171), .Y(n2237) );
  OAI2BB2X2 U864 ( .B0(n2040), .B1(n264), .A0N(n2040), .A1N(n2039), .Y(n2054)
         );
  NAND3X1 U865 ( .A(n316), .B(n1948), .C(n2446), .Y(n2040) );
  NAND2X1 U866 ( .A(n744), .B(n367), .Y(n607) );
  INVXL U867 ( .A(n2231), .Y(n165) );
  CLKINVX1 U868 ( .A(n165), .Y(n166) );
  NOR2BX1 U869 ( .AN(n2405), .B(n2399), .Y(n2409) );
  OAI2BB2X2 U870 ( .B0(n2393), .B1(work_cntr[15]), .A0N(n2393), .A1N(
        work_cntr[15]), .Y(n2399) );
  OAI22X2 U871 ( .A0(n2488), .A1(n2487), .B0(n2486), .B1(n2485), .Y(n2494) );
  OAI21X1 U872 ( .A0(n2465), .A1(n264), .B0(n2464), .Y(n2480) );
  NAND2X1 U873 ( .A(n2465), .B(n264), .Y(n2464) );
  OAI21X2 U874 ( .A0(n1977), .A1(n1976), .B0(n1981), .Y(n1992) );
  NAND2X1 U875 ( .A(n1976), .B(n1968), .Y(n1981) );
  CLKINVX1 U876 ( .A(n927), .Y(n923) );
  CLKINVX1 U877 ( .A(n167), .Y(n168) );
  CLKINVX1 U878 ( .A(n2637), .Y(n2636) );
  AOI21X1 U879 ( .A0(n270), .A1(n1008), .B0(n1007), .Y(n2637) );
  OAI31X4 U880 ( .A0(n2286), .A1(n2309), .A2(n2285), .B0(n2284), .Y(n2334) );
  CLKINVX1 U881 ( .A(n2310), .Y(n2285) );
  OAI2BB2X1 U882 ( .B0(write_addr[13]), .B1(n1811), .A0N(write_addr[13]), 
        .A1N(n1811), .Y(n2766) );
  NOR2X2 U883 ( .A(n235), .B(n2820), .Y(n1811) );
  AND2X2 U884 ( .A(n371), .B(n370), .Y(n603) );
  NAND2X1 U885 ( .A(n744), .B(n368), .Y(n371) );
  OAI21X1 U886 ( .A0(n2715), .A1(n2711), .B0(write_addr[9]), .Y(n2714) );
  NAND2BX1 U887 ( .AN(n2854), .B(n2715), .Y(n2755) );
  NOR2X1 U888 ( .A(n2715), .B(n317), .Y(n2708) );
  NOR2X2 U889 ( .A(n235), .B(n1825), .Y(n2715) );
  CLKINVX1 U890 ( .A(n845), .Y(n826) );
  OAI31X1 U891 ( .A0(n1325), .A1(n1324), .A2(n1323), .B0(n1322), .Y(n1333) );
  OAI21X2 U892 ( .A0(n1313), .A1(n2423), .B0(n1312), .Y(n1324) );
  CLKINVX1 U893 ( .A(n2000), .Y(n169) );
  CLKINVX1 U894 ( .A(n2575), .Y(n2571) );
  OAI21X1 U895 ( .A0(n1002), .A1(work_cntr[11]), .B0(n1001), .Y(n2575) );
  AND2X2 U896 ( .A(n2085), .B(n2084), .Y(n2099) );
  NOR2BX2 U897 ( .AN(n2125), .B(n2124), .Y(n2149) );
  NOR2X1 U898 ( .A(n2165), .B(n2121), .Y(n2125) );
  NAND2X1 U899 ( .A(curr_photo_size[1]), .B(curr_photo_size[0]), .Y(n2867) );
  AOI2BB2X2 U900 ( .B0(n1079), .B1(n1078), .A0N(n1079), .A1N(n1078), .Y(n1124)
         );
  NAND2X1 U901 ( .A(n1042), .B(n1034), .Y(n1079) );
  OAI31X1 U902 ( .A0(n1048), .A1(n1047), .A2(n227), .B0(n1050), .Y(n1062) );
  NAND2X1 U903 ( .A(n1047), .B(n227), .Y(n1050) );
  NAND3X1 U904 ( .A(n744), .B(n366), .C(n365), .Y(n619) );
  NOR2X2 U905 ( .A(n1214), .B(n1216), .Y(n1270) );
  NOR2X2 U906 ( .A(N1827), .B(n1193), .Y(n1214) );
  OAI2BB2X2 U907 ( .B0(work_cntr[14]), .B1(n1312), .A0N(work_cntr[14]), .A1N(
        n1312), .Y(n1316) );
  NAND2X1 U908 ( .A(n1313), .B(n2423), .Y(n1312) );
  OAI31X4 U909 ( .A0(n1301), .A1(n1297), .A2(n1300), .B0(n1295), .Y(n1306) );
  OAI21X2 U910 ( .A0(n1294), .A1(n1293), .B0(n1296), .Y(n1300) );
  OAI21X1 U911 ( .A0(n1966), .A1(n2128), .B0(n1965), .Y(n1976) );
  NOR2X1 U912 ( .A(n1965), .B(next_work_cntr[16]), .Y(n1959) );
  OAI2BB2X2 U913 ( .B0(next_work_cntr[16]), .B1(n1965), .A0N(
        next_work_cntr[16]), .A1N(n1965), .Y(n1971) );
  NAND2X1 U914 ( .A(n2128), .B(n1966), .Y(n1965) );
  NOR2BX1 U915 ( .AN(n967), .B(n966), .Y(n969) );
  NOR2X2 U916 ( .A(n962), .B(n965), .Y(n966) );
  CLKINVX1 U917 ( .A(n962), .Y(n1802) );
  OAI21X1 U918 ( .A0(n960), .A1(n262), .B0(n947), .Y(n962) );
  CLKINVX1 U919 ( .A(n1923), .Y(n170) );
  OAI22X1 U920 ( .A0(n1363), .A1(n1362), .B0(n1361), .B1(n1360), .Y(n1368) );
  OAI22X2 U921 ( .A0(n1340), .A1(n266), .B0(n1354), .B1(n2380), .Y(n1362) );
  NOR2BX2 U922 ( .AN(n1567), .B(n1566), .Y(n1588) );
  NAND2X1 U923 ( .A(write_cntr[9]), .B(n277), .Y(n1567) );
  NOR2X1 U924 ( .A(write_cntr[9]), .B(n277), .Y(n1566) );
  OAI22X2 U925 ( .A0(write_cntr[0]), .A1(n961), .B0(n220), .B1(n960), .Y(n1892) );
  NAND2X1 U926 ( .A(n316), .B(n961), .Y(n960) );
  AOI2BB2X2 U927 ( .B0(n1142), .B1(n1141), .A0N(n1142), .A1N(n1141), .Y(n1168)
         );
  NAND2BX1 U928 ( .AN(n1110), .B(n1109), .Y(n1142) );
  CLKINVX1 U929 ( .A(n2620), .Y(n2619) );
  OAI21X1 U930 ( .A0(n1713), .A1(n261), .B0(n1709), .Y(n1714) );
  CLKINVX1 U931 ( .A(n1713), .Y(n2380) );
  NAND2X2 U932 ( .A(n1713), .B(n261), .Y(n1709) );
  NOR2X2 U933 ( .A(work_cntr[8]), .B(n1723), .Y(n1713) );
  NOR2X2 U934 ( .A(n317), .B(n2520), .Y(next_work_cntr[17]) );
  OAI22X1 U935 ( .A0(n2519), .A1(n2518), .B0(n2520), .B1(n259), .Y(n2531) );
  CLKINVX1 U936 ( .A(n2519), .Y(n2520) );
  CLKINVX1 U937 ( .A(n2601), .Y(n2600) );
  AOI21X1 U938 ( .A0(n1005), .A1(n266), .B0(n1004), .Y(n2601) );
  AOI21X1 U939 ( .A0(work_cntr[18]), .A1(n2379), .B0(n1643), .Y(n1653) );
  OAI21X2 U940 ( .A0(n1643), .A1(n259), .B0(n1788), .Y(n1651) );
  NAND2BX1 U941 ( .AN(n1169), .B(n1161), .Y(n1196) );
  NAND2X1 U942 ( .A(n1160), .B(n1189), .Y(n1169) );
  INVXL U943 ( .A(n1115), .Y(n171) );
  CLKINVX1 U944 ( .A(n171), .Y(n172) );
  NOR2X1 U945 ( .A(n1191), .B(n1192), .Y(n1185) );
  NAND2BX1 U946 ( .AN(n1172), .B(n1170), .Y(n1191) );
  OAI21X2 U947 ( .A0(n1646), .A1(n257), .B0(n1645), .Y(n1650) );
  NAND2X1 U948 ( .A(write_addr[9]), .B(write_addr[10]), .Y(n2854) );
  OAI21X1 U949 ( .A0(n2119), .A1(n2522), .B0(next_work_cntr[18]), .Y(n2134) );
  NAND2BX1 U950 ( .AN(next_work_cntr[18]), .B(n1960), .Y(n1958) );
  NOR2X2 U951 ( .A(n317), .B(n2521), .Y(next_work_cntr[18]) );
  OAI211X1 U952 ( .A0(work_cntr[19]), .A1(n231), .B0(n257), .C0(n1407), .Y(
        n1414) );
  AOI31X1 U953 ( .A0(work_cntr[18]), .A1(n1407), .A2(n1414), .B0(n1413), .Y(
        n1410) );
  NAND2X1 U954 ( .A(n2518), .B(n231), .Y(n1407) );
  NAND2X1 U955 ( .A(n2476), .B(n2382), .Y(n2393) );
  CLKINVX1 U956 ( .A(n1877), .Y(n1805) );
  OAI22X1 U957 ( .A0(n1877), .A1(n933), .B0(n932), .B1(n931), .Y(n948) );
  OAI22X1 U958 ( .A0(n1805), .A1(n2754), .B0(n1877), .B1(n2761), .Y(n944) );
  AOI221X4 U959 ( .A0(n276), .A1(n929), .B0(n317), .B1(n929), .C0(n834), .Y(
        n1877) );
  AOI2BB2X2 U960 ( .B0(n1956), .B1(n1746), .A0N(n1956), .A1N(n1746), .Y(n1759)
         );
  NOR2BX1 U961 ( .AN(n1956), .B(n1746), .Y(n1753) );
  NOR2X2 U962 ( .A(n317), .B(n1956), .Y(n2060) );
  OAI21X2 U963 ( .A0(n270), .A1(n221), .B0(n2446), .Y(n1956) );
  OAI2BB2X2 U964 ( .B0(n2044), .B1(n2042), .A0N(n2044), .A1N(n2042), .Y(n2065)
         );
  OAI31X4 U965 ( .A0(n2719), .A1(n241), .A2(n855), .B0(n854), .Y(n861) );
  OAI22X1 U966 ( .A0(n1807), .A1(n2719), .B0(n1018), .B1(n2720), .Y(n869) );
  NAND2X1 U967 ( .A(n2718), .B(n2719), .Y(n2723) );
  CLKINVX1 U968 ( .A(n2720), .Y(n2719) );
  NOR2BX1 U969 ( .AN(n1969), .B(next_work_cntr[14]), .Y(n1966) );
  NOR2X2 U970 ( .A(n317), .B(n2545), .Y(next_work_cntr[14]) );
  CLKINVX1 U971 ( .A(n2582), .Y(n2581) );
  AOI21X2 U972 ( .A0(n1003), .A1(n228), .B0(n1002), .Y(n2582) );
  OAI22X2 U973 ( .A0(work_cntr[4]), .A1(n2476), .B0(n270), .B1(n2477), .Y(
        n2495) );
  NOR2X2 U974 ( .A(n2378), .B(N1827), .Y(n2476) );
  NOR2X2 U975 ( .A(n2664), .B(n317), .Y(next_work_cntr[1]) );
  NOR4BX1 U976 ( .AN(n2313), .B(next_work_cntr[1]), .C(n2329), .D(n2328), .Y(
        n2337) );
  NOR2X1 U977 ( .A(next_work_cntr[1]), .B(n2340), .Y(n2372) );
  CLKINVX1 U978 ( .A(n877), .Y(n1804) );
  NOR2X2 U979 ( .A(n317), .B(n2658), .Y(next_work_cntr[2]) );
  CLKINVX1 U980 ( .A(\DP_OP_229J1_126_7015/I3 ), .Y(n173) );
  OA21X2 U981 ( .A0(n2493), .A1(n2503), .B0(n2492), .Y(n2506) );
  OAI221X4 U982 ( .A0(n2503), .A1(n2502), .B0(n2501), .B1(n2500), .C0(n2499), 
        .Y(n2507) );
  OAI21X2 U983 ( .A0(n273), .A1(n2496), .B0(n2477), .Y(n2503) );
  CLKINVX1 U984 ( .A(n2137), .Y(next_work_cntr[8]) );
  NAND2X1 U985 ( .A(n2027), .B(n2137), .Y(n2018) );
  OAI2BB2X1 U986 ( .B0(n2137), .B1(n2027), .A0N(n2137), .A1N(n2027), .Y(n2035)
         );
  NAND2X2 U987 ( .A(n316), .B(n2601), .Y(n2137) );
  OAI21X1 U988 ( .A0(n1644), .A1(n231), .B0(n2379), .Y(n1665) );
  NAND2X2 U989 ( .A(n1644), .B(n231), .Y(n2379) );
  NOR2X1 U990 ( .A(next_work_cntr[19]), .B(n1958), .Y(n2109) );
  NAND2BX1 U991 ( .AN(n2114), .B(next_work_cntr[19]), .Y(n2115) );
  OAI2BB2X2 U992 ( .B0(next_work_cntr[19]), .B1(n1958), .A0N(
        next_work_cntr[19]), .A1N(n1958), .Y(n1972) );
  NOR2X2 U993 ( .A(n317), .B(n2522), .Y(next_work_cntr[19]) );
  AOI32X4 U994 ( .A0(n1972), .A1(n1964), .A2(n1963), .B0(n1971), .B1(n1964), 
        .Y(n1982) );
  CLKINVX1 U995 ( .A(n1855), .Y(n1873) );
  OAI22X2 U996 ( .A0(write_cntr[5]), .A1(n836), .B0(n274), .B1(n835), .Y(n1855) );
  OAI22X1 U997 ( .A0(n2722), .A1(n1015), .B0(n2724), .B1(n1806), .Y(n874) );
  NOR2X1 U998 ( .A(n1806), .B(n1938), .Y(n1016) );
  OAI22X2 U999 ( .A0(n1015), .A1(n1938), .B0(n1806), .B1(next_cr_x[6]), .Y(
        n1832) );
  CLKINVX1 U1000 ( .A(n1015), .Y(n1806) );
  NAND2X1 U1001 ( .A(n2145), .B(n2153), .Y(n2124) );
  NAND2X2 U1002 ( .A(n316), .B(n2563), .Y(n2153) );
  NAND2X1 U1003 ( .A(write_addr[16]), .B(n369), .Y(n370) );
  AND2X2 U1004 ( .A(n27), .B(n748), .Y(n747) );
  OAI21X1 U1005 ( .A0(n27), .A1(n2111), .B0(n789), .Y(n799) );
  NAND2X1 U1006 ( .A(n27), .B(n798), .Y(n803) );
  AND2X2 U1007 ( .A(n27), .B(en_so), .Y(n742) );
  NOR2X2 U1008 ( .A(n317), .B(n2526), .Y(next_work_cntr[16]) );
  NAND2X2 U1009 ( .A(n1020), .B(n1019), .Y(next_cr_x[5]) );
  NOR2X1 U1010 ( .A(n1925), .B(n1929), .Y(n1940) );
  CLKINVX1 U1011 ( .A(n1926), .Y(n1929) );
  AOI2BB2X2 U1012 ( .B0(n829), .B1(n828), .A0N(n829), .A1N(n828), .Y(n1014) );
  OAI22X1 U1013 ( .A0(n2718), .A1(n844), .B0(n226), .B1(n829), .Y(n852) );
  INVX3 U1014 ( .A(n844), .Y(n829) );
  AOI2BB2X2 U1015 ( .B0(next_work_cntr[7]), .B1(n1957), .A0N(next_work_cntr[7]), .A1N(n1957), .Y(n2044) );
  NOR2X1 U1016 ( .A(next_work_cntr[7]), .B(n1957), .Y(n2027) );
  NOR2X2 U1017 ( .A(n317), .B(n2613), .Y(next_work_cntr[7]) );
  INVX3 U1018 ( .A(\next_cr_y[0] ), .Y(n174) );
  OR2X2 U1019 ( .A(n727), .B(n726), .Y(n728) );
  OR2X2 U1020 ( .A(n2853), .B(\sftr_n[0]_BAR ), .Y(n717) );
  NAND2X1 U1021 ( .A(n266), .B(n1085), .Y(n1100) );
  NOR2X1 U1022 ( .A(n266), .B(n1085), .Y(n1101) );
  BUFX4 U1023 ( .A(n133), .Y(n315) );
  CLKINVX1 U1024 ( .A(n2145), .Y(next_work_cntr[11]) );
  NAND2X1 U1025 ( .A(write_addr[8]), .B(n2848), .Y(n1808) );
  NAND2X1 U1026 ( .A(write_addr[8]), .B(n2831), .Y(n1813) );
  NOR2X1 U1027 ( .A(n2847), .B(write_addr[8]), .Y(n2843) );
  NAND2X2 U1028 ( .A(n221), .B(n270), .Y(n2446) );
  NOR2X1 U1029 ( .A(n221), .B(n1143), .Y(n1172) );
  OAI22X2 U1030 ( .A0(n1280), .A1(n221), .B0(n1354), .B1(n2446), .Y(n1386) );
  INVX3 U1031 ( .A(n1783), .Y(n724) );
  OAI211X4 U1032 ( .A0(n1393), .A1(n2654), .B0(n1392), .C0(n1391), .Y(n1405)
         );
  NOR2X2 U1033 ( .A(n317), .B(n2654), .Y(next_work_cntr[3]) );
  NAND2X2 U1034 ( .A(n1008), .B(n1354), .Y(n2654) );
  OAI21X4 U1035 ( .A0(write_cntr[4]), .A1(n834), .B0(n835), .Y(n1880) );
  NOR2X1 U1036 ( .A(n836), .B(n317), .Y(n835) );
  OAI21X1 U1037 ( .A0(n2783), .A1(n2681), .B0(n2682), .Y(n946) );
  AOI2BB2X2 U1038 ( .B0(n310), .B1(\intadd_3/SUM[6] ), .A0N(n2783), .A1N(n364), 
        .Y(n650) );
  INVX3 U1039 ( .A(n744), .Y(n2783) );
  INVX16 U1040 ( .A(n8), .Y(cr_a[2]) );
  INVX16 U1041 ( .A(n4), .Y(cr_a[0]) );
  CLKINVX1 U1042 ( .A(n2883), .Y(n177) );
  INVX16 U1043 ( .A(n177), .Y(cr_a[3]) );
  OAI22X2 U1044 ( .A0(work_cntr[4]), .A1(n1354), .B0(n270), .B1(n1402), .Y(
        n1387) );
  INVX16 U1045 ( .A(n6), .Y(cr_a[1]) );
  CLKINVX1 U1046 ( .A(n2882), .Y(n180) );
  INVX16 U1047 ( .A(n180), .Y(cr_a[4]) );
  CLKINVX1 U1048 ( .A(n2881), .Y(n182) );
  INVX16 U1049 ( .A(n182), .Y(cr_a[5]) );
  CLKINVX1 U1050 ( .A(n2880), .Y(n184) );
  INVX16 U1051 ( .A(n184), .Y(cr_a[6]) );
  CLKINVX1 U1052 ( .A(n2879), .Y(n186) );
  INVX16 U1053 ( .A(n186), .Y(cr_a[7]) );
  INVX16 U1054 ( .A(n9), .Y(cr_a[8]) );
  OAI22X1 U1055 ( .A0(n216), .A1(n1046), .B0(work_cntr[14]), .B1(n1035), .Y(
        n1061) );
  NOR2X1 U1056 ( .A(work_cntr[14]), .B(n1072), .Y(n1047) );
  OAI2BB2X1 U1057 ( .B0(n1072), .B1(work_cntr[14]), .A0N(n1072), .A1N(n1071), 
        .Y(n1106) );
  NAND2X1 U1058 ( .A(n998), .B(work_cntr[14]), .Y(n997) );
  AND2X2 U1059 ( .A(n747), .B(n379), .Y(n740) );
  INVX3 U1060 ( .A(n652), .Y(n718) );
  NOR2X2 U1061 ( .A(read_cntr[0]), .B(n286), .Y(n652) );
  CLKINVX1 U1062 ( .A(n2878), .Y(n189) );
  INVX16 U1063 ( .A(n189), .Y(im_wen_n) );
  AOI31XL U1064 ( .A0(n1796), .A1(n306), .A2(n1795), .B0(n1794), .Y(n2878) );
  NAND2X1 U1065 ( .A(write_addr[12]), .B(n2762), .Y(n2765) );
  NOR2X1 U1066 ( .A(n2756), .B(n2755), .Y(n2762) );
  AND2XL U1067 ( .A(n531), .B(n774), .Y(n420) );
  CLKINVX1 U1068 ( .A(n420), .Y(n191) );
  OAI31X4 U1069 ( .A0(n419), .A1(n774), .A2(n418), .B0(n191), .Y(n512) );
  AOI21X1 U1070 ( .A0(n2695), .A1(n2686), .B0(n2694), .Y(n2685) );
  CLKINVX1 U1071 ( .A(n2690), .Y(n2694) );
  NAND2BX1 U1072 ( .AN(n1209), .B(n1212), .Y(n1213) );
  NAND2BX1 U1073 ( .AN(n1495), .B(n1497), .Y(n1501) );
  NOR2X1 U1074 ( .A(n1489), .B(n1494), .Y(n1495) );
  NAND2X1 U1075 ( .A(n1261), .B(n1230), .Y(n1236) );
  NOR2BX1 U1076 ( .AN(n2768), .B(n2773), .Y(n2769) );
  NOR2X1 U1077 ( .A(work_cntr[4]), .B(n1164), .Y(n1189) );
  NOR2BX1 U1078 ( .AN(n1166), .B(n1165), .Y(n1164) );
  AOI211X1 U1079 ( .A0(n248), .A1(n323), .B0(n324), .C0(n783), .Y(n760) );
  NAND2X1 U1080 ( .A(global_cntr[13]), .B(n322), .Y(n323) );
  NAND2X1 U1081 ( .A(n2180), .B(n2179), .Y(n2207) );
  OAI21X1 U1082 ( .A0(n1528), .A1(n1527), .B0(n263), .Y(n1533) );
  NOR2BX1 U1083 ( .AN(n1534), .B(n1528), .Y(n1536) );
  NOR2X1 U1084 ( .A(n1526), .B(n1525), .Y(n1528) );
  NOR2X1 U1085 ( .A(n225), .B(cr_read_cntr[7]), .Y(n1023) );
  OAI21X1 U1086 ( .A0(n2670), .A1(n2665), .B0(n2664), .Y(n2667) );
  NOR2X1 U1087 ( .A(n2666), .B(n2665), .Y(n2669) );
  NOR2BX1 U1088 ( .AN(n2663), .B(n2662), .Y(n2665) );
  CLKINVX1 U1089 ( .A(n1593), .Y(n1609) );
  OAI21X1 U1090 ( .A0(n1648), .A1(n1649), .B0(n1650), .Y(n1663) );
  OAI21X2 U1091 ( .A0(n1649), .A1(n1650), .B0(n1663), .Y(n1676) );
  NOR2X1 U1092 ( .A(n1657), .B(n1647), .Y(n1649) );
  NOR2X1 U1093 ( .A(n1715), .B(n1714), .Y(n1724) );
  NAND2X1 U1094 ( .A(n994), .B(work_cntr[18]), .Y(n2516) );
  OAI21X2 U1095 ( .A0(n994), .A1(work_cntr[18]), .B0(n2516), .Y(n2521) );
  NOR2X1 U1096 ( .A(n995), .B(n231), .Y(n994) );
  NOR2X1 U1097 ( .A(n1659), .B(n1658), .Y(n1664) );
  NOR2X1 U1098 ( .A(n2699), .B(n2696), .Y(n2697) );
  NAND2X1 U1099 ( .A(n2692), .B(cr_read_cntr[5]), .Y(n2696) );
  NOR2BX1 U1100 ( .AN(n1758), .B(n1759), .Y(n1751) );
  NOR2X1 U1101 ( .A(work_cntr[4]), .B(n1749), .Y(n1758) );
  NOR2X1 U1102 ( .A(n278), .B(n819), .Y(n816) );
  AOI211X1 U1103 ( .A0(n278), .A1(n819), .B0(n816), .C0(n317), .Y(n844) );
  NAND3X1 U1104 ( .A(write_cntr[9]), .B(write_cntr[10]), .C(n821), .Y(n819) );
  NOR2BX1 U1105 ( .AN(n2831), .B(n2853), .Y(n2833) );
  OAI31X1 U1106 ( .A0(n1132), .A1(n1158), .A2(n1128), .B0(n1137), .Y(n1135) );
  NAND2BX1 U1107 ( .AN(n1130), .B(n1129), .Y(n1158) );
  NOR2BX1 U1108 ( .AN(n1843), .B(n1937), .Y(n1844) );
  NOR2X1 U1109 ( .A(n1685), .B(n1684), .Y(n1694) );
  OAI21X1 U1110 ( .A0(n1682), .A1(n1681), .B0(n1680), .Y(n1684) );
  NOR4X1 U1111 ( .A(n2329), .B(n2353), .C(n2356), .D(next_work_cntr[0]), .Y(
        n2361) );
  OAI2BB2X1 U1112 ( .B0(n2330), .B1(n2331), .A0N(n2330), .A1N(n2328), .Y(n2356) );
  OAI21X1 U1113 ( .A0(n2253), .A1(n2252), .B0(n2251), .Y(n2271) );
  OAI21X1 U1114 ( .A0(n1488), .A1(n1487), .B0(n1486), .Y(n1494) );
  OAI21X1 U1115 ( .A0(n268), .A1(n1483), .B0(n1487), .Y(n1492) );
  OAI21X1 U1116 ( .A0(n1482), .A1(n1481), .B0(n268), .Y(n1487) );
  OAI222X4 U1117 ( .A0(n238), .A1(n2771), .B0(n776), .B1(n2834), .C0(n1917), 
        .C1(n1916), .Y(n713) );
  OAI21X1 U1118 ( .A0(write_addr[2]), .A1(write_addr[1]), .B0(n1915), .Y(n2834) );
  OAI21X1 U1119 ( .A0(n2711), .A1(n2843), .B0(n1825), .Y(n2707) );
  OAI211X1 U1120 ( .A0(n2782), .A1(n1821), .B0(n1820), .C0(n1819), .Y(n1825)
         );
  OAI21X1 U1121 ( .A0(n2822), .A1(n2853), .B0(n2851), .Y(n2821) );
  NAND2X2 U1122 ( .A(n2795), .B(n2842), .Y(n2853) );
  NAND2X2 U1123 ( .A(n316), .B(n1947), .Y(n2771) );
  NOR2XL U1124 ( .A(n807), .B(n1947), .Y(n745) );
  NOR2X2 U1125 ( .A(next_state[2]), .B(next_state[1]), .Y(n1947) );
  OAI211X1 U1126 ( .A0(n538), .A1(n555), .B0(n537), .C0(n536), .Y(\C1/Z_1 ) );
  CLKINVX1 U1127 ( .A(n2170), .Y(n2203) );
  NOR2X1 U1128 ( .A(n2170), .B(n2200), .Y(n2183) );
  OAI22X1 U1129 ( .A0(n2137), .A1(n2136), .B0(next_work_cntr[8]), .B1(n2143), 
        .Y(n2170) );
  NOR2XL U1130 ( .A(n2662), .B(n2657), .Y(n193) );
  OAI21X2 U1131 ( .A0(n2658), .A1(n2663), .B0(n192), .Y(n2672) );
  NOR2X1 U1132 ( .A(n2656), .B(n2655), .Y(n2662) );
  OAI21X4 U1133 ( .A0(N1826), .A1(n1789), .B0(n1397), .Y(n2658) );
  OAI21X1 U1134 ( .A0(n1229), .A1(n1228), .B0(n1227), .Y(n1230) );
  OAI22X1 U1135 ( .A0(n1207), .A1(n1206), .B0(n1205), .B1(n1204), .Y(n1228) );
  OAI21X1 U1136 ( .A0(n2274), .A1(n2273), .B0(n2272), .Y(n2303) );
  OAI21X1 U1137 ( .A0(n2291), .A1(n2249), .B0(n2273), .Y(n2272) );
  OAI22X1 U1138 ( .A0(n2248), .A1(n2247), .B0(n2250), .B1(n2246), .Y(n2273) );
  AOI22X2 U1139 ( .A0(n1261), .A1(n1260), .B0(n1264), .B1(n1259), .Y(n1551) );
  OAI22X1 U1140 ( .A0(n1243), .A1(n1274), .B0(n1242), .B1(n1241), .Y(n1264) );
  OAI22X1 U1141 ( .A0(n2083), .A1(n2082), .B0(n2081), .B1(n2080), .Y(n2084) );
  OAI22X1 U1142 ( .A0(n2080), .A1(n2073), .B0(n2072), .B1(n2071), .Y(n2076) );
  OAI22X1 U1143 ( .A0(n2074), .A1(n2071), .B0(n2075), .B1(n2069), .Y(n2080) );
  OAI2BB2X1 U1144 ( .B0(n1065), .B1(n1064), .A0N(n1065), .A1N(n1064), .Y(n1094) );
  OAI21X1 U1145 ( .A0(n1739), .A1(n1736), .B0(n1735), .Y(n1747) );
  NOR2X1 U1146 ( .A(n1736), .B(n1735), .Y(n1741) );
  OAI2BB2X1 U1147 ( .B0(n1570), .B1(n1569), .A0N(n1570), .A1N(n1569), .Y(n1579) );
  NAND3X1 U1148 ( .A(n1570), .B(n1565), .C(n1562), .Y(n1572) );
  AOI2BB2X2 U1149 ( .B0(write_cntr[11]), .B1(n1559), .A0N(write_cntr[11]), 
        .A1N(n1559), .Y(n1570) );
  NOR2X1 U1150 ( .A(n1642), .B(n1036), .Y(n1035) );
  NAND2X1 U1151 ( .A(n507), .B(n468), .Y(n508) );
  XOR2X1 U1152 ( .A(n526), .B(curr_time[18]), .Y(n507) );
  MXI2X1 U1153 ( .A(n538), .B(n399), .S0(curr_time[10]), .Y(n503) );
  OA21X1 U1154 ( .A0(n400), .A1(n398), .B0(n405), .Y(n538) );
  AOI2BB2X2 U1155 ( .B0(n251), .B1(n1081), .A0N(n251), .A1N(n1081), .Y(n1084)
         );
  OAI21X2 U1156 ( .A0(n1043), .A1(n1044), .B0(n1042), .Y(n1081) );
  NAND2X1 U1157 ( .A(n1558), .B(n277), .Y(n1560) );
  AND2X2 U1158 ( .A(write_cntr[14]), .B(n1561), .Y(n277) );
  AOI22X1 U1159 ( .A0(work_cntr[11]), .A1(n1327), .B0(n1402), .B1(n2414), .Y(
        n1336) );
  CLKINVX1 U1160 ( .A(n1689), .Y(n2414) );
  CLKINVX1 U1161 ( .A(n710), .Y(n696) );
  OR2X4 U1162 ( .A(n569), .B(n719), .Y(n710) );
  NAND2X1 U1163 ( .A(n2875), .B(n2874), .Y(so_mux_sel[0]) );
  OAI2BB2X1 U1164 ( .B0(curr_time[12]), .B1(m_1[3]), .A0N(curr_time[12]), 
        .A1N(m_1[3]), .Y(n983) );
  NAND2X1 U1165 ( .A(n341), .B(n345), .Y(m_1[3]) );
  AOI21X1 U1166 ( .A0(n243), .A1(n327), .B0(n328), .Y(n754) );
  NAND2X1 U1167 ( .A(n392), .B(n395), .Y(m_1[2]) );
  NOR2X1 U1168 ( .A(n347), .B(n346), .Y(n395) );
  AOI2BB2X2 U1169 ( .B0(n1592), .B1(n1591), .A0N(n1592), .A1N(n1591), .Y(n1611) );
  NOR3X1 U1170 ( .A(n287), .B(n1592), .C(n1593), .Y(n1595) );
  NAND2BX1 U1171 ( .AN(n1586), .B(n1584), .Y(n1592) );
  NOR2X1 U1172 ( .A(n739), .B(n738), .Y(n2810) );
  NOR2X1 U1173 ( .A(n384), .B(n2864), .Y(n739) );
  NOR2X1 U1174 ( .A(n1594), .B(n287), .Y(n1605) );
  NOR2X1 U1175 ( .A(n1691), .B(n1690), .Y(n1699) );
  NAND2X1 U1176 ( .A(n546), .B(n1800), .Y(n553) );
  NAND2X1 U1177 ( .A(n743), .B(n546), .Y(n554) );
  NOR2X1 U1178 ( .A(n424), .B(n1801), .Y(n546) );
  OAI22X1 U1179 ( .A0(n414), .A1(n989), .B0(n990), .B1(n991), .Y(n418) );
  NOR2X1 U1180 ( .A(n355), .B(n354), .Y(n414) );
  NOR2X1 U1181 ( .A(n1138), .B(n1170), .Y(n1149) );
  NAND2X1 U1182 ( .A(n221), .B(n1143), .Y(n1170) );
  NOR2X1 U1183 ( .A(n2089), .B(n2098), .Y(n2091) );
  CLKINVX1 U1184 ( .A(n2087), .Y(n2098) );
  OAI2BB2X1 U1185 ( .B0(n1182), .B1(n1181), .A0N(n1182), .A1N(n1181), .Y(n1207) );
  NOR2BX1 U1186 ( .AN(n1182), .B(n1181), .Y(n1184) );
  NOR2BX1 U1187 ( .AN(n1178), .B(n1177), .Y(n1181) );
  NOR2BX1 U1188 ( .AN(n1266), .B(n1268), .Y(n1279) );
  NAND2X1 U1189 ( .A(n263), .B(n1212), .Y(n1266) );
  NOR2X1 U1190 ( .A(n263), .B(n1212), .Y(n1268) );
  NOR2X1 U1191 ( .A(n1375), .B(n1374), .Y(n1383) );
  OAI21X1 U1192 ( .A0(n1375), .A1(n1371), .B0(n1370), .Y(n1374) );
  NOR2BX1 U1193 ( .AN(n2155), .B(n2157), .Y(n2191) );
  NOR2X1 U1194 ( .A(n2236), .B(n2233), .Y(n2239) );
  CLKINVX1 U1195 ( .A(n1931), .Y(n776) );
  AOI211X4 U1196 ( .A0(n1931), .A1(\next_write_addr_w[0] ), .B0(n1895), .C0(
        n376), .Y(n716) );
  NOR2X1 U1197 ( .A(n1823), .B(n1944), .Y(n1931) );
  NOR2X1 U1198 ( .A(next_work_cntr[13]), .B(n1985), .Y(n1969) );
  CLKINVX1 U1199 ( .A(n2116), .Y(next_work_cntr[13]) );
  NOR2X1 U1200 ( .A(n1892), .B(n1900), .Y(n1908) );
  NAND2X1 U1201 ( .A(n1006), .B(work_cntr[7]), .Y(n1005) );
  OAI21X2 U1202 ( .A0(n1006), .A1(work_cntr[7]), .B0(n1005), .Y(n2613) );
  AOI21X1 U1203 ( .A0(n1948), .A1(n264), .B0(n1006), .Y(n2620) );
  NOR2X1 U1204 ( .A(n1948), .B(n264), .Y(n1006) );
  NOR2X1 U1205 ( .A(n2406), .B(n2405), .Y(n2418) );
  NAND2X1 U1206 ( .A(n996), .B(work_cntr[16]), .Y(n995) );
  OAI21X2 U1207 ( .A0(n996), .A1(work_cntr[16]), .B0(n995), .Y(n2526) );
  NOR2X1 U1208 ( .A(n997), .B(n227), .Y(n996) );
  OAI21X1 U1209 ( .A0(n2860), .A1(n2859), .B0(n2873), .Y(n2871) );
  NOR2X1 U1210 ( .A(n1772), .B(n263), .Y(n2860) );
  NOR2X1 U1211 ( .A(n2477), .B(n2446), .Y(n2465) );
  CLKINVX1 U1212 ( .A(n2476), .Y(n2477) );
  OAI2BB2X1 U1213 ( .B0(n2029), .B1(n2028), .A0N(n2029), .A1N(n2028), .Y(n2049) );
  NOR2BX1 U1214 ( .AN(n2029), .B(n2028), .Y(n2031) );
  OAI2BB2X1 U1215 ( .B0(n2025), .B1(n2024), .A0N(n2025), .A1N(n2023), .Y(n2029) );
  AOI21X2 U1216 ( .A0(n1933), .A1(n1804), .B0(n1829), .Y(n1850) );
  NOR2X1 U1217 ( .A(n1804), .B(n1933), .Y(n1829) );
  NAND2BX1 U1218 ( .AN(next_work_cntr[10]), .B(n2009), .Y(n1998) );
  NOR2X1 U1219 ( .A(n136), .B(n2018), .Y(n2009) );
  NOR2X1 U1220 ( .A(n1988), .B(n1987), .Y(n2001) );
  AOI2BB2X2 U1221 ( .B0(next_work_cntr[2]), .B1(n2305), .A0N(next_work_cntr[2]), .A1N(n2305), .Y(n2371) );
  NOR2X1 U1222 ( .A(next_work_cntr[2]), .B(n2305), .Y(n2312) );
  NOR2BX1 U1223 ( .AN(n2323), .B(n2324), .Y(n2305) );
  AOI21X1 U1224 ( .A0(work_cntr[8]), .A1(n1723), .B0(n1713), .Y(n1726) );
  NOR2X1 U1225 ( .A(n1555), .B(n1640), .Y(N2292) );
  NAND2X1 U1226 ( .A(global_cntr[2]), .B(n1554), .Y(n1640) );
  OAI21X1 U1227 ( .A0(curr_time[15]), .A1(n772), .B0(n977), .Y(n979) );
  NOR2X1 U1228 ( .A(n259), .B(n1401), .Y(n1413) );
  OAI21X1 U1229 ( .A0(curr_time[23]), .A1(n771), .B0(n971), .Y(n973) );
  AND2X2 U1230 ( .A(global_cntr[1]), .B(global_cntr[0]), .Y(n769) );
  NOR3X1 U1231 ( .A(global_cntr[1]), .B(n253), .C(n1640), .Y(N2272) );
  NAND2X1 U1232 ( .A(global_cntr[1]), .B(n253), .Y(n1555) );
  NOR4X2 U1233 ( .A(global_cntr[0]), .B(global_cntr[1]), .C(n1640), .D(N2294), 
        .Y(en_photo_num) );
  OAI21X1 U1234 ( .A0(n2387), .A1(n252), .B0(n2386), .Y(n2390) );
  NAND2X1 U1235 ( .A(n2387), .B(n252), .Y(n2386) );
  NOR2X1 U1236 ( .A(n2477), .B(n2379), .Y(n2387) );
  OAI21X1 U1237 ( .A0(n2481), .A1(n2480), .B0(n2479), .Y(n2486) );
  OAI2BB2X1 U1238 ( .B0(n2469), .B1(n2468), .A0N(n2469), .A1N(n2467), .Y(n2481) );
  OAI21X1 U1239 ( .A0(n2788), .A1(n2787), .B0(n2786), .Y(n2793) );
  AOI22X1 U1240 ( .A0(n310), .A1(\intadd_3/SUM[7] ), .B0(n2716), .B1(n2755), 
        .Y(n2850) );
  OA21X2 U1241 ( .A0(n463), .A1(n466), .B0(n460), .Y(n526) );
  OAI21X1 U1242 ( .A0(n459), .A1(n460), .B0(n467), .Y(n471) );
  OAI21X1 U1243 ( .A0(n1359), .A1(n1362), .B0(n1369), .Y(n1366) );
  OAI2BB2X1 U1244 ( .B0(n1350), .B1(n1349), .A0N(n1350), .A1N(n1348), .Y(n1359) );
  AOI2BB2X2 U1245 ( .B0(n310), .B1(\intadd_3/SUM[0] ), .A0N(n776), .A1N(n2835), 
        .Y(n701) );
  OAI21X1 U1246 ( .A0(n1986), .A1(n2153), .B0(n1985), .Y(n1997) );
  NOR2X1 U1247 ( .A(next_work_cntr[11]), .B(n1998), .Y(n1986) );
  NAND2X1 U1248 ( .A(n1986), .B(n2153), .Y(n1985) );
  NAND2BX1 U1249 ( .AN(n2059), .B(n2063), .Y(n2072) );
  OAI21X1 U1250 ( .A0(n2056), .A1(n2055), .B0(n2054), .Y(n2063) );
  OAI31X1 U1251 ( .A0(n1437), .A1(work_cntr[13]), .A2(n1436), .B0(n1435), .Y(
        n1444) );
  OAI21X1 U1252 ( .A0(n216), .A1(n1430), .B0(n1429), .Y(n1436) );
  OAI31X4 U1253 ( .A0(n2629), .A1(n2628), .A2(n2627), .B0(n2626), .Y(n2635) );
  OAI21X1 U1254 ( .A0(n2619), .A1(n2618), .B0(n2623), .Y(n2627) );
  OAI21X1 U1255 ( .A0(n2600), .A1(n2599), .B0(n2604), .Y(n2608) );
  OAI22X1 U1256 ( .A0(n852), .A1(n851), .B0(n857), .B1(n850), .Y(n864) );
  OAI21X1 U1257 ( .A0(n219), .A1(n849), .B0(n848), .Y(n857) );
  OAI21X1 U1258 ( .A0(n1028), .A1(n1027), .B0(cr_read_cntr[4]), .Y(n1032) );
  OAI21X1 U1259 ( .A0(n2581), .A1(n2580), .B0(n2585), .Y(n2589) );
  OAI21X1 U1260 ( .A0(n217), .A1(n1447), .B0(n1446), .Y(n1452) );
  OAI21X1 U1261 ( .A0(n2562), .A1(n2561), .B0(n2566), .Y(n2570) );
  OAI21X1 U1262 ( .A0(curr_time[18]), .A1(n526), .B0(n462), .Y(n467) );
  NOR2X1 U1263 ( .A(n462), .B(curr_time[18]), .Y(n466) );
  OAI21X1 U1264 ( .A0(n974), .A1(n513), .B0(n455), .Y(n462) );
  NOR2X1 U1265 ( .A(n1908), .B(n1907), .Y(n1905) );
  AOI22X1 U1266 ( .A0(n967), .A1(n966), .B0(n965), .B1(n964), .Y(n1907) );
  CLKINVX1 U1267 ( .A(n1692), .Y(n1704) );
  OAI21X1 U1268 ( .A0(n1695), .A1(n1690), .B0(n1691), .Y(n1692) );
  OAI21X1 U1269 ( .A0(n2198), .A1(n2196), .B0(n2194), .Y(n2219) );
  OAI21X1 U1270 ( .A0(n2163), .A1(n2162), .B0(n2161), .Y(n2198) );
  NOR2X1 U1271 ( .A(n2781), .B(n2780), .Y(n2784) );
  AOI211X4 U1272 ( .A0(n2781), .A1(n2780), .B0(n2784), .C0(n2783), .Y(n2830)
         );
  OAI21X1 U1273 ( .A0(write_addr[18]), .A1(n1814), .B0(n1813), .Y(n2781) );
  OAI21X1 U1274 ( .A0(n1316), .A1(n1314), .B0(n1309), .Y(n1321) );
  OAI22X1 U1275 ( .A0(n1306), .A1(n1305), .B0(n1304), .B1(n1308), .Y(n1314) );
  OAI22X1 U1276 ( .A0(n155), .A1(n1617), .B0(n1613), .B1(n1612), .Y(n1637) );
  CLKINVX1 U1277 ( .A(n2174), .Y(n2172) );
  NOR2X1 U1278 ( .A(n2174), .B(n2164), .Y(n2154) );
  NOR2BX1 U1279 ( .AN(n2175), .B(n2174), .Y(n2211) );
  OAI22X1 U1280 ( .A0(n2145), .A1(n2144), .B0(next_work_cntr[11]), .B1(n2123), 
        .Y(n2174) );
  AOI22X1 U1281 ( .A0(n1618), .A1(n1617), .B0(n1616), .B1(n155), .Y(n1638) );
  OAI22X1 U1282 ( .A0(n1598), .A1(n1597), .B0(n1601), .B1(n1596), .Y(n1618) );
  OAI22X1 U1283 ( .A0(n2199), .A1(n2198), .B0(n2197), .B1(n2196), .Y(n2220) );
  OAI22X1 U1284 ( .A0(n2193), .A1(n2142), .B0(n2141), .B1(n2160), .Y(n2199) );
  OAI22X1 U1285 ( .A0(n223), .A1(n1808), .B0(write_addr[11]), .B1(n2713), .Y(
        n2756) );
  NAND3X1 U1286 ( .A(n1720), .B(n1710), .C(n1716), .Y(n1712) );
  AOI2BB2X2 U1287 ( .B0(n1707), .B1(n1706), .A0N(n1707), .A1N(n1706), .Y(n1720) );
  MXI2X2 U1288 ( .A(n397), .B(n400), .S0(n396), .Y(n533) );
  NOR2X1 U1289 ( .A(n401), .B(curr_time[10]), .Y(n400) );
  NOR2X1 U1290 ( .A(n2317), .B(n2316), .Y(n2341) );
  NOR2X2 U1291 ( .A(n942), .B(n949), .Y(n2717) );
  MXI2X2 U1292 ( .A(n987), .B(curr_time[3]), .S0(n988), .Y(n992) );
  AND2X2 U1293 ( .A(n413), .B(n414), .Y(n988) );
  AOI211X4 U1294 ( .A0(n240), .A1(n330), .B0(n329), .C0(n783), .Y(n753) );
  NOR2X2 U1295 ( .A(n782), .B(n781), .Y(n783) );
  NOR2X2 U1296 ( .A(n194), .B(n195), .Y(n1946) );
  OAI21X1 U1297 ( .A0(n254), .A1(n1555), .B0(n1946), .Y(n801) );
  NAND2X1 U1298 ( .A(n767), .B(n1946), .Y(n2111) );
  NAND4BX1 U1299 ( .AN(n768), .B(n1947), .C(n1946), .D(n1945), .Y(n2790) );
  AOI211X4 U1300 ( .A0(n218), .A1(n334), .B0(n336), .C0(n783), .Y(n750) );
  AOI211X4 U1301 ( .A0(n250), .A1(n325), .B0(n758), .C0(n783), .Y(n757) );
  AOI2BB2X2 U1302 ( .B0(n466), .B1(n976), .A0N(n465), .A1N(n464), .Y(n520) );
  NAND2BX1 U1303 ( .AN(n2261), .B(n2260), .Y(n2309) );
  NAND2X1 U1304 ( .A(n142), .B(n2223), .Y(n2260) );
  NAND2X1 U1305 ( .A(n268), .B(n1092), .Y(n1109) );
  NOR2X1 U1306 ( .A(n2012), .B(n2013), .Y(n2025) );
  NAND2BX1 U1307 ( .AN(n2013), .B(n2019), .Y(n2033) );
  NOR2X2 U1308 ( .A(n2008), .B(n2007), .Y(n2013) );
  OAI21X1 U1309 ( .A0(n2006), .A1(n2005), .B0(n2004), .Y(n2007) );
  NAND2BX1 U1310 ( .AN(next_work_cntr[7]), .B(n2180), .Y(n2200) );
  NOR2BX1 U1311 ( .AN(next_work_cntr[7]), .B(n2180), .Y(n2201) );
  OAI2BB2X1 U1312 ( .B0(n1108), .B1(n1107), .A0N(n1108), .A1N(n1107), .Y(n1137) );
  NOR2X2 U1313 ( .A(n1063), .B(n1062), .Y(n1108) );
  NOR2X2 U1314 ( .A(n232), .B(n263), .Y(n2378) );
  NOR2BX2 U1315 ( .AN(n416), .B(n415), .Y(n524) );
  NOR2X2 U1316 ( .A(n1798), .B(write_cntr[5]), .Y(n1629) );
  BUFX2 U1317 ( .A(n1693), .Y(n196) );
  NOR3BX1 U1318 ( .AN(n196), .B(n1688), .C(n1702), .Y(n1695) );
  INVXL U1319 ( .A(n1568), .Y(n198) );
  NOR2X1 U1320 ( .A(n198), .B(n199), .Y(n200) );
  NOR2XL U1321 ( .A(write_cntr[10]), .B(n1568), .Y(n201) );
  OAI2BB2X1 U1322 ( .B0(n197), .B1(n1582), .A0N(n197), .A1N(n1582), .Y(n1598)
         );
  NAND3X1 U1323 ( .A(n1577), .B(n197), .C(n1579), .Y(n1580) );
  NOR2BX2 U1324 ( .AN(n2032), .B(n2026), .Y(n2030) );
  NAND2X1 U1325 ( .A(n2021), .B(n2020), .Y(n2032) );
  NOR2X1 U1326 ( .A(n2021), .B(n2020), .Y(n2026) );
  NOR2BX2 U1327 ( .AN(n2135), .B(n2133), .Y(n2165) );
  NAND2X1 U1328 ( .A(n316), .B(n2590), .Y(n2120) );
  NAND2X1 U1329 ( .A(n202), .B(n203), .Y(n1148) );
  INVXL U1330 ( .A(n1111), .Y(n204) );
  INVXL U1331 ( .A(n1112), .Y(n205) );
  NAND2XL U1332 ( .A(n1112), .B(n1111), .Y(n202) );
  NAND2X1 U1333 ( .A(n204), .B(n205), .Y(n203) );
  OAI2BB2X1 U1334 ( .B0(n1149), .B1(n1148), .A0N(n1149), .A1N(n1148), .Y(n1197) );
  NAND2X1 U1335 ( .A(n1149), .B(n1148), .Y(n1179) );
  NAND2BX1 U1336 ( .AN(n1101), .B(n1100), .Y(n1112) );
  OAI21X1 U1337 ( .A0(n1110), .A1(n1139), .B0(n1109), .Y(n1111) );
  AOI211X1 U1338 ( .A0(n1771), .A1(n1770), .B0(n1769), .C0(n318), .Y(
        expand_sel[1]) );
  NOR2BX2 U1339 ( .AN(n2122), .B(n2124), .Y(n2146) );
  AOI2BB2X2 U1340 ( .B0(n2116), .B1(n2146), .A0N(n2116), .A1N(n2146), .Y(n2155) );
  NAND2X1 U1341 ( .A(n206), .B(n207), .Y(n2335) );
  CLKINVX1 U1342 ( .A(n2281), .Y(n208) );
  INVXL U1343 ( .A(n2282), .Y(n209) );
  NAND2XL U1344 ( .A(n2282), .B(n2281), .Y(n206) );
  NAND2X1 U1345 ( .A(n208), .B(n209), .Y(n207) );
  NOR2X1 U1346 ( .A(n2335), .B(n2366), .Y(n2313) );
  NOR2BX1 U1347 ( .AN(n2336), .B(n2335), .Y(n2316) );
  CLKINVX1 U1348 ( .A(n2289), .Y(n2282) );
  CLKINVX1 U1349 ( .A(n210), .Y(n2319) );
  NOR2X1 U1350 ( .A(n2319), .B(n2318), .Y(n2297) );
  AOI2BB2X2 U1351 ( .B0(n2238), .B1(n2239), .A0N(n2238), .A1N(n2239), .Y(n2291) );
  OA21X1 U1352 ( .A0(n2594), .A1(n2595), .B0(n2593), .Y(n2605) );
  CLKINVX1 U1353 ( .A(n2594), .Y(n2590) );
  OAI21X2 U1354 ( .A0(n1004), .A1(work_cntr[9]), .B0(n1003), .Y(n2594) );
  NAND2X1 U1355 ( .A(n1004), .B(work_cntr[9]), .Y(n1003) );
  OAI2BB2X2 U1356 ( .B0(n1848), .B1(n1925), .A0N(n1848), .A1N(n1925), .Y(n1859) );
  AO21X2 U1357 ( .A0(n272), .A1(n839), .B0(n838), .Y(n1848) );
  NOR2XL U1358 ( .A(n1730), .B(n268), .Y(n213) );
  INVXL U1359 ( .A(n1723), .Y(n214) );
  NAND2X1 U1360 ( .A(n1730), .B(n268), .Y(n1723) );
  OAI2BB2X1 U1361 ( .B0(n1233), .B1(n1232), .A0N(n1233), .A1N(n1232), .Y(n1247) );
  NAND2BX1 U1362 ( .AN(n1232), .B(n1233), .Y(n1210) );
  NAND2X1 U1363 ( .A(n1233), .B(n1245), .Y(n1244) );
  AOI2BB2X2 U1364 ( .B0(n1169), .B1(n1168), .A0N(n1169), .A1N(n1168), .Y(n1233) );
  AOI2BB2X2 U1365 ( .B0(n2265), .B1(n2264), .A0N(n2265), .A1N(n2264), .Y(n2307) );
  AOI2BB2X2 U1366 ( .B0(n1200), .B1(n1199), .A0N(n1200), .A1N(n1198), .Y(n1241) );
  OAI2BB2X1 U1367 ( .B0(n1199), .B1(n1179), .A0N(n1199), .A1N(n1179), .Y(n1198) );
  NOR2X1 U1368 ( .A(n1199), .B(n1156), .Y(n1152) );
  NOR2X1 U1369 ( .A(n1199), .B(n1179), .Y(n1153) );
  NOR2X1 U1370 ( .A(n1199), .B(n1196), .Y(n1176) );
  AOI2BB2X2 U1371 ( .B0(n172), .B1(n1114), .A0N(n172), .A1N(n1114), .Y(n1199)
         );
  OAI21X2 U1372 ( .A0(n1074), .A1(n1073), .B0(n1105), .Y(n1132) );
  NOR2XL U1373 ( .A(n1846), .B(n1937), .Y(n215) );
  CLKINVX1 U1374 ( .A(n1941), .Y(n1937) );
  NOR3X1 U1375 ( .A(n1855), .B(n131), .C(n1859), .Y(n1866) );
  CLKINVX1 U1376 ( .A(n1846), .Y(n1857) );
  NAND2X2 U1377 ( .A(n1852), .B(n1851), .Y(n1941) );
  OAI211X4 U1378 ( .A0(write_cntr[6]), .A1(n837), .B0(n316), .C0(n839), .Y(
        n1846) );
  CLKINVX1 U1379 ( .A(n2664), .Y(n2668) );
  CLKINVX1 U1380 ( .A(n1807), .Y(n1018) );
  NAND2X1 U1381 ( .A(n819), .B(n818), .Y(n1807) );
  CLKINVX1 U1382 ( .A(n2383), .Y(n1283) );
  NOR2BX2 U1383 ( .AN(n930), .B(n812), .Y(n837) );
  NAND2X1 U1384 ( .A(write_cntr[2]), .B(n930), .Y(n929) );
  OAI211X4 U1385 ( .A0(write_cntr[2]), .A1(n930), .B0(n316), .C0(n929), .Y(
        n1803) );
  NOR3X2 U1386 ( .A(n262), .B(n220), .C(n961), .Y(n930) );
  CLKINVX1 U1387 ( .A(n946), .Y(n961) );
  NAND2X2 U1388 ( .A(n316), .B(n2535), .Y(n2128) );
  AOI21X2 U1389 ( .A0(n997), .A1(n227), .B0(n996), .Y(n2535) );
  NAND2X1 U1390 ( .A(n2827), .B(write_addr[17]), .Y(n2829) );
  NOR3X2 U1391 ( .A(n2820), .B(n2824), .C(n280), .Y(n2827) );
  NAND2X1 U1392 ( .A(write_addr[13]), .B(n2774), .Y(n2824) );
  CLKINVX1 U1393 ( .A(n2748), .Y(n2744) );
  NAND2X1 U1394 ( .A(n908), .B(n910), .Y(n2748) );
  CLKINVX1 U1395 ( .A(n2737), .Y(n2742) );
  NAND2X1 U1396 ( .A(n902), .B(n2737), .Y(n906) );
  NAND2X2 U1397 ( .A(n903), .B(n898), .Y(n2737) );
  AOI21X1 U1398 ( .A0(n1830), .A1(n2704), .B0(n1829), .Y(n1831) );
  CLKINVX1 U1399 ( .A(n2704), .Y(n1925) );
  NAND2X2 U1400 ( .A(n1837), .B(n1836), .Y(n2704) );
  OAI31X4 U1401 ( .A0(n2241), .A1(n2243), .A2(n2242), .B0(n2240), .Y(n2298) );
  NOR2BX1 U1402 ( .AN(n2239), .B(n2238), .Y(n2242) );
  NOR3X1 U1403 ( .A(n1112), .B(n1142), .C(work_cntr[6]), .Y(n1113) );
  NOR2X2 U1404 ( .A(work_cntr[6]), .B(n2446), .Y(n1730) );
  NOR2X2 U1405 ( .A(work_cntr[10]), .B(n1709), .Y(n1705) );
  OAI21X1 U1406 ( .A0(n1705), .A1(n251), .B0(n1689), .Y(n1707) );
  OAI2BB2X1 U1407 ( .B0(n1328), .B1(n228), .A0N(n1402), .A1N(n1705), .Y(n1338)
         );
  NAND2X1 U1408 ( .A(n1705), .B(n251), .Y(n1689) );
  CLKINVX1 U1409 ( .A(n2724), .Y(n2722) );
  NOR2X2 U1410 ( .A(n862), .B(n861), .Y(n2724) );
  CLKINVX1 U1411 ( .A(n2733), .Y(n2730) );
  OAI22X1 U1412 ( .A0(n2735), .A1(n2734), .B0(n2733), .B1(n2732), .Y(n2741) );
  NOR2X2 U1413 ( .A(n888), .B(n887), .Y(n2733) );
  NAND2X1 U1414 ( .A(n2212), .B(n2210), .Y(n2214) );
  OAI2BB2X2 U1415 ( .B0(n2213), .B1(n2212), .A0N(n2213), .A1N(n2212), .Y(n2245) );
  NOR2X2 U1416 ( .A(n2190), .B(n2178), .Y(n2212) );
  NOR2X1 U1417 ( .A(n2154), .B(n2148), .Y(n2178) );
  AND2X2 U1418 ( .A(n2154), .B(n2153), .Y(n2190) );
  NOR2X2 U1419 ( .A(n1800), .B(n549), .Y(n552) );
  NOR2X1 U1420 ( .A(n1222), .B(n1198), .Y(n1203) );
  NOR2X1 U1421 ( .A(n1222), .B(n1244), .Y(n1240) );
  OAI21X2 U1422 ( .A0(n1163), .A1(n1162), .B0(n1196), .Y(n1222) );
  OAI2BB2X1 U1423 ( .B0(n1237), .B1(n1213), .A0N(n1237), .A1N(n1213), .Y(n1253) );
  OAI21X1 U1424 ( .A0(n1237), .A1(n1208), .B0(n1228), .Y(n1227) );
  NOR2X1 U1425 ( .A(n1237), .B(n1213), .Y(n1234) );
  OAI2BB2X2 U1426 ( .B0(n1191), .B1(n1190), .A0N(n1191), .A1N(n1190), .Y(n1237) );
  OAI21X1 U1427 ( .A0(n1189), .A1(n1214), .B0(n1188), .Y(n1190) );
  OAI2BB2X1 U1428 ( .B0(n2728), .B1(n2727), .A0N(n2728), .A1N(n2727), .Y(n2732) );
  CLKINVX1 U1429 ( .A(n2728), .Y(n2725) );
  NAND2X2 U1430 ( .A(n873), .B(n883), .Y(n2728) );
  NOR2X2 U1431 ( .A(n2855), .B(n2854), .Y(n2848) );
  OAI21X1 U1432 ( .A0(n1817), .A1(write_addr[7]), .B0(n2855), .Y(n2840) );
  CLKINVX1 U1433 ( .A(n2855), .Y(n2847) );
  NOR2X1 U1434 ( .A(n2855), .B(n235), .Y(n2711) );
  NAND2X2 U1435 ( .A(n1817), .B(write_addr[7]), .Y(n2855) );
  CLKINVX1 U1436 ( .A(n1788), .Y(n1771) );
  AND2X2 U1437 ( .A(n566), .B(n565), .Y(n725) );
  NAND2XL U1438 ( .A(n1786), .B(n740), .Y(n566) );
  OAI31X4 U1439 ( .A0(n2278), .A1(n2277), .A2(n2295), .B0(n2276), .Y(n2343) );
  NOR2X1 U1440 ( .A(n2761), .B(n2760), .Y(n2759) );
  CLKINVX1 U1441 ( .A(n2761), .Y(n2754) );
  NOR2X2 U1442 ( .A(n928), .B(n163), .Y(n2761) );
  NOR2X2 U1443 ( .A(\sftr_n[0]_BAR ), .B(n2851), .Y(n707) );
  CLKINVX1 U1444 ( .A(n2841), .Y(n2851) );
  CLKINVX1 U1445 ( .A(n1936), .Y(n1932) );
  OAI21X2 U1446 ( .A0(n1909), .A1(n1936), .B0(n1927), .Y(n1924) );
  NAND2X2 U1447 ( .A(n1870), .B(n1869), .Y(n1936) );
  NAND3X1 U1448 ( .A(N196), .B(n2378), .C(N1827), .Y(n1008) );
  NOR2X1 U1449 ( .A(N1825), .B(N196), .Y(n1772) );
  AOI221X4 U1450 ( .A0(n1771), .A1(N196), .B0(n1775), .B1(n284), .C0(n318), 
        .Y(expand_sel[0]) );
  OAI22X1 U1451 ( .A0(N196), .A1(n1551), .B0(n284), .B1(n1278), .Y(n2863) );
  OAI21X2 U1452 ( .A0(n2035), .A1(n2034), .B0(n2036), .Y(n2057) );
  NOR2BX1 U1453 ( .AN(n2037), .B(n2048), .Y(n2036) );
  CLKINVX1 U1454 ( .A(n2128), .Y(next_work_cntr[15]) );
  NAND2X1 U1455 ( .A(n922), .B(n2752), .Y(n925) );
  OAI21X1 U1456 ( .A0(n2750), .A1(n2752), .B0(n2749), .Y(n2758) );
  NAND2X2 U1457 ( .A(n917), .B(n918), .Y(n2752) );
  INVX3 U1458 ( .A(n723), .Y(n700) );
  AND2X2 U1459 ( .A(n581), .B(n740), .Y(n723) );
  OAI22X2 U1460 ( .A0(n1000), .A1(work_cntr[12]), .B0(n1001), .B1(n217), .Y(
        n2562) );
  OAI22X1 U1461 ( .A0(work_cntr[12]), .A1(n2414), .B0(n217), .B1(n1689), .Y(
        n1688) );
  CLKINVX1 U1462 ( .A(next_cr_x[6]), .Y(n1938) );
  OAI22X1 U1463 ( .A0(n1016), .A1(n1829), .B0(n1015), .B1(next_cr_x[6]), .Y(
        n1017) );
  CLKINVX2 U1464 ( .A(n831), .Y(next_cr_x[6]) );
  NOR2X2 U1465 ( .A(n2855), .B(n236), .Y(n2804) );
  CLKINVX1 U1466 ( .A(n2695), .Y(n2699) );
  NOR2BX4 U1467 ( .AN(next_en_si), .B(n2682), .Y(n2695) );
  NAND2BX1 U1468 ( .AN(n1928), .B(n1896), .Y(n1910) );
  AOI22X4 U1469 ( .A0(n1891), .A1(n1890), .B0(n1889), .B1(n1888), .Y(n1928) );
  CLKINVX2 U1470 ( .A(n715), .Y(n697) );
  NAND2BX2 U1471 ( .AN(curr_photo_size[0]), .B(read_cntr[0]), .Y(n715) );
  AOI211X4 U1472 ( .A0(write_cntr[9]), .A1(n821), .B0(n317), .C0(n820), .Y(
        n1015) );
  INVX6 U1473 ( .A(n2086), .Y(n317) );
  NAND2X4 U1474 ( .A(n569), .B(n737), .Y(n704) );
  NAND2X4 U1475 ( .A(n273), .B(n1397), .Y(n1354) );
  NAND2X1 U1476 ( .A(N1826), .B(n1789), .Y(n1397) );
  AND2X4 U1477 ( .A(n2857), .B(n740), .Y(n720) );
  AND2X4 U1478 ( .A(n1783), .B(n339), .Y(n746) );
  NOR2X2 U1479 ( .A(n1555), .B(n1639), .Y(N2250) );
  NAND2X1 U1480 ( .A(n1554), .B(n254), .Y(n1639) );
  NAND3X2 U1481 ( .A(n27), .B(n26), .C(n229), .Y(N2294) );
  NAND2XL U1482 ( .A(curr_photo[0]), .B(n304), .Y(n381) );
  NOR2XL U1483 ( .A(curr_photo[0]), .B(n2793), .Y(n2791) );
  NOR2XL U1484 ( .A(n2789), .B(n2790), .Y(n2786) );
  NOR2BX1 U1485 ( .AN(N1141), .B(n318), .Y(n2883) );
  NOR2BXL U1486 ( .AN(N1142), .B(n318), .Y(n2882) );
  NOR2BXL U1487 ( .AN(N1143), .B(n318), .Y(n2881) );
  NOR2BXL U1488 ( .AN(N1144), .B(n318), .Y(n2880) );
  NOR2BXL U1489 ( .AN(N1145), .B(n318), .Y(n2879) );
  NAND4XL U1490 ( .A(n496), .B(n484), .C(n483), .D(n474), .Y(\C1/Z_3 ) );
  NAND2XL U1491 ( .A(n532), .B(\s_1[3] ), .Y(n474) );
  OAI211XL U1492 ( .A0(n508), .A1(n471), .B0(n552), .C0(n470), .Y(n483) );
  INVXL U1493 ( .A(n541), .Y(n469) );
  INVXL U1494 ( .A(n466), .Y(n459) );
  AOI22XL U1495 ( .A0(n551), .A1(n425), .B0(n550), .B1(n426), .Y(n484) );
  XOR2XL U1496 ( .A(n423), .B(n422), .Y(n425) );
  NOR2XL U1497 ( .A(n545), .B(n510), .Y(n423) );
  XNOR2XL U1498 ( .A(n407), .B(n406), .Y(n408) );
  OAI211XL U1499 ( .A0(n405), .A1(n404), .B0(n403), .C0(n402), .Y(n406) );
  NAND2XL U1500 ( .A(n538), .B(n401), .Y(n402) );
  INVXL U1501 ( .A(n400), .Y(n404) );
  NOR2XL U1502 ( .A(n539), .B(n501), .Y(n407) );
  AOI21XL U1503 ( .A0(n552), .A1(n517), .B0(n516), .Y(n518) );
  INVXL U1504 ( .A(n513), .Y(n514) );
  AOI22XL U1505 ( .A0(n512), .A1(n511), .B0(n524), .B1(n510), .Y(n515) );
  NAND2XL U1506 ( .A(n524), .B(n509), .Y(n511) );
  INVXL U1507 ( .A(curr_time[1]), .Y(n509) );
  NOR2XL U1508 ( .A(n520), .B(curr_time[17]), .Y(n506) );
  AOI22XL U1509 ( .A0(n505), .A1(m_1[2]), .B0(n540), .B1(n504), .Y(n519) );
  NAND2XL U1510 ( .A(n405), .B(n398), .Y(n399) );
  INVXL U1511 ( .A(n555), .Y(n505) );
  OAI211XL U1512 ( .A0(n539), .A1(n535), .B0(n540), .C0(n534), .Y(n536) );
  NAND2XL U1513 ( .A(n533), .B(n535), .Y(n534) );
  INVXL U1514 ( .A(curr_time[9]), .Y(n535) );
  AOI211XL U1515 ( .A0(n532), .A1(n531), .B0(n530), .C0(n529), .Y(n537) );
  INVXL U1516 ( .A(n550), .Y(n525) );
  MXI2XL U1517 ( .A(n524), .B(n545), .S0(curr_time[1]), .Y(n527) );
  INVXL U1518 ( .A(n551), .Y(n528) );
  AOI211XL U1519 ( .A0(curr_time[17]), .A1(n541), .B0(n523), .C0(n522), .Y(
        n530) );
  NOR2XL U1520 ( .A(curr_time[17]), .B(n521), .Y(n522) );
  INVXL U1521 ( .A(n520), .Y(n521) );
  INVXL U1522 ( .A(n552), .Y(n523) );
  INVXL U1523 ( .A(n553), .Y(n532) );
  INVXL U1524 ( .A(n562), .Y(n559) );
  NOR3XL U1525 ( .A(n552), .B(n551), .C(n550), .Y(n556) );
  AOI21XL U1526 ( .A0(n552), .A1(\h_0[0] ), .B0(n542), .Y(n543) );
  INVXL U1527 ( .A(n463), .Y(n464) );
  AOI21XL U1528 ( .A0(n462), .A1(curr_time[18]), .B0(n461), .Y(n465) );
  INVXL U1529 ( .A(n460), .Y(n461) );
  NAND2XL U1530 ( .A(n513), .B(n974), .Y(n455) );
  INVXL U1531 ( .A(curr_time[19]), .Y(n974) );
  INVXL U1532 ( .A(n431), .Y(n432) );
  NOR2XL U1533 ( .A(n430), .B(n429), .Y(n433) );
  INVXL U1534 ( .A(curr_time[22]), .Y(n429) );
  NAND2XL U1535 ( .A(n975), .B(n428), .Y(n458) );
  NOR2XL U1536 ( .A(curr_time[21]), .B(curr_time[22]), .Y(n972) );
  NAND2BXL U1537 ( .AN(n973), .B(n427), .Y(n430) );
  INVXL U1538 ( .A(curr_time[20]), .Y(n427) );
  NAND3XL U1539 ( .A(curr_time[23]), .B(curr_time[22]), .C(n771), .Y(n971) );
  INVXL U1540 ( .A(curr_time[21]), .Y(n771) );
  INVXL U1541 ( .A(curr_time[17]), .Y(n468) );
  NAND2XL U1542 ( .A(n1800), .B(n409), .Y(n548) );
  INVXL U1543 ( .A(n1801), .Y(n409) );
  INVXL U1544 ( .A(n424), .Y(n410) );
  NAND2XL U1545 ( .A(n1622), .B(n1799), .Y(n1797) );
  NAND2XL U1546 ( .A(n403), .B(n405), .Y(n397) );
  NAND2XL U1547 ( .A(n401), .B(curr_time[10]), .Y(n403) );
  INVXL U1548 ( .A(n396), .Y(n398) );
  NAND2XL U1549 ( .A(n389), .B(n388), .Y(n390) );
  INVXL U1550 ( .A(n982), .Y(n388) );
  INVXL U1551 ( .A(n395), .Y(n389) );
  INVXL U1552 ( .A(n983), .Y(n391) );
  INVXL U1553 ( .A(n981), .Y(n386) );
  NAND2XL U1554 ( .A(n980), .B(m_1[2]), .Y(n981) );
  NOR2XL U1555 ( .A(m_1[2]), .B(n980), .Y(n387) );
  INVXL U1556 ( .A(n345), .Y(n346) );
  NOR2XL U1557 ( .A(n344), .B(n343), .Y(n347) );
  INVXL U1558 ( .A(curr_time[14]), .Y(n343) );
  NAND2XL U1559 ( .A(n983), .B(n980), .Y(n982) );
  INVXL U1560 ( .A(curr_time[11]), .Y(n980) );
  NOR2XL U1561 ( .A(curr_time[13]), .B(curr_time[14]), .Y(n978) );
  NAND3XL U1562 ( .A(n344), .B(curr_time[14]), .C(n340), .Y(n341) );
  NAND2BXL U1563 ( .AN(curr_time[13]), .B(curr_time[15]), .Y(n340) );
  NAND2BXL U1564 ( .AN(n979), .B(n342), .Y(n344) );
  INVXL U1565 ( .A(curr_time[12]), .Y(n342) );
  NAND3XL U1566 ( .A(curr_time[15]), .B(curr_time[14]), .C(n772), .Y(n977) );
  INVXL U1567 ( .A(curr_time[13]), .Y(n772) );
  NAND2XL U1568 ( .A(n1799), .B(n1798), .Y(n1801) );
  AOI211XL U1569 ( .A0(n1635), .A1(n1634), .B0(n1633), .C0(n1632), .Y(n1636)
         );
  INVXL U1570 ( .A(n1618), .Y(n1616) );
  INVXL U1571 ( .A(n1637), .Y(n1614) );
  NAND2BXL U1572 ( .AN(n1607), .B(n1606), .Y(n1608) );
  AND2XL U1573 ( .A(n1624), .B(n1637), .Y(n1635) );
  NOR2XL U1574 ( .A(n1611), .B(n1610), .Y(n1612) );
  NAND4BXL U1575 ( .AN(n1629), .B(write_cntr[4]), .C(n1607), .D(n1606), .Y(
        n1624) );
  INVXL U1576 ( .A(n1798), .Y(n1622) );
  INVXL U1577 ( .A(n1585), .Y(n1590) );
  NOR2XL U1578 ( .A(n1600), .B(n1599), .Y(n1597) );
  INVXL U1579 ( .A(n1594), .Y(n1619) );
  INVXL U1580 ( .A(n1602), .Y(n1596) );
  NOR2BXL U1581 ( .AN(n197), .B(n1582), .Y(n1578) );
  INVXL U1582 ( .A(n1576), .Y(n1581) );
  NAND2XL U1583 ( .A(n1585), .B(n1589), .Y(n1593) );
  NAND2XL U1584 ( .A(n1583), .B(n272), .Y(n1589) );
  AND2XL U1585 ( .A(n1575), .B(n1580), .Y(n1574) );
  NOR2BXL U1586 ( .AN(n1570), .B(n1569), .Y(n1564) );
  INVXL U1587 ( .A(n1571), .Y(n1563) );
  AOI211XL U1588 ( .A0(curr_time[2]), .A1(n417), .B0(n419), .C0(n418), .Y(n415) );
  NAND2XL U1589 ( .A(n421), .B(n416), .Y(n531) );
  NAND2XL U1590 ( .A(n418), .B(n993), .Y(n416) );
  NAND2XL U1591 ( .A(n992), .B(n774), .Y(n993) );
  INVXL U1592 ( .A(curr_time[2]), .Y(n774) );
  NOR2XL U1593 ( .A(curr_time[3]), .B(n988), .Y(n990) );
  INVXL U1594 ( .A(n419), .Y(n421) );
  NAND2XL U1595 ( .A(n411), .B(n414), .Y(n412) );
  INVXL U1596 ( .A(n992), .Y(n417) );
  INVXL U1597 ( .A(n353), .Y(n354) );
  NOR2XL U1598 ( .A(n352), .B(n351), .Y(n355) );
  INVXL U1599 ( .A(curr_time[6]), .Y(n351) );
  NAND2XL U1600 ( .A(n991), .B(n987), .Y(n989) );
  NOR2XL U1601 ( .A(curr_time[5]), .B(curr_time[6]), .Y(n985) );
  NAND3XL U1602 ( .A(n352), .B(curr_time[6]), .C(n348), .Y(n349) );
  NAND2BXL U1603 ( .AN(curr_time[5]), .B(curr_time[7]), .Y(n348) );
  NAND2BXL U1604 ( .AN(n986), .B(n350), .Y(n352) );
  INVXL U1605 ( .A(curr_time[4]), .Y(n350) );
  NAND3XL U1606 ( .A(curr_time[7]), .B(curr_time[6]), .C(n773), .Y(n984) );
  INVXL U1607 ( .A(curr_time[5]), .Y(n773) );
  INVXL U1608 ( .A(curr_time[3]), .Y(n987) );
  NOR2XL U1609 ( .A(n1033), .B(n302), .Y(n558) );
  MXI2XL U1610 ( .A(cr_read_cntr[4]), .B(n1032), .S0(n1033), .Y(n563) );
  INVXL U1611 ( .A(n1029), .Y(n1031) );
  INVXL U1612 ( .A(n561), .Y(n564) );
  NAND2XL U1613 ( .A(n560), .B(cr_read_cntr[3]), .Y(n561) );
  NAND2XL U1614 ( .A(n1032), .B(n557), .Y(n560) );
  NAND2XL U1615 ( .A(n1030), .B(n1029), .Y(n1027) );
  NAND2XL U1616 ( .A(cr_read_cntr[5]), .B(n1026), .Y(n1029) );
  NOR3XL U1617 ( .A(cr_read_cntr[7]), .B(n301), .C(n225), .Y(n1025) );
  INVXL U1618 ( .A(n1023), .Y(n1024) );
  AOI22XL U1619 ( .A0(n1781), .A1(n1780), .B0(n1792), .B1(n1788), .Y(n1782) );
  NOR2XL U1620 ( .A(n273), .B(n1775), .Y(n1781) );
  NOR2BXL U1621 ( .AN(n1780), .B(n2860), .Y(n1773) );
  INVXL U1622 ( .A(n1790), .Y(n1769) );
  NAND2XL U1623 ( .A(n2664), .B(n1951), .Y(n1770) );
  OAI211XL U1624 ( .A0(n2873), .A1(n2872), .B0(n737), .C0(n2871), .Y(n2874) );
  NAND3XL U1625 ( .A(n740), .B(n2864), .C(n2863), .Y(n2865) );
  INVXL U1626 ( .A(n2862), .Y(n2866) );
  NOR4XL U1627 ( .A(n2861), .B(n263), .C(n2867), .D(n2871), .Y(n2870) );
  MXI2XL U1628 ( .A(n2877), .B(n2876), .S0(read_cntr[0]), .Y(n473) );
  NAND3XL U1629 ( .A(next_en_si), .B(n744), .C(n306), .Y(n2877) );
  OAI211XL U1630 ( .A0(n2687), .A1(cr_read_cntr[3]), .B0(n2695), .C0(n2689), 
        .Y(n2688) );
  OAI211XL U1631 ( .A0(n2692), .A1(cr_read_cntr[5]), .B0(n2695), .C0(n2696), 
        .Y(n2693) );
  NOR2XL U1632 ( .A(n2685), .B(n380), .Y(n453) );
  NAND2X1 U1633 ( .A(N1139), .B(N1138), .Y(n2686) );
  INVXL U1634 ( .A(n2702), .Y(n2700) );
  NAND2XL U1635 ( .A(cr_read_cntr[6]), .B(n2697), .Y(n2702) );
  AOI211XL U1636 ( .A0(n2678), .A1(n740), .B0(n2677), .C0(n2676), .Y(n2679) );
  NAND2XL U1637 ( .A(n2660), .B(n192), .Y(n2659) );
  INVXL U1638 ( .A(n2661), .Y(n2657) );
  NOR2XL U1639 ( .A(n138), .B(n2660), .Y(n2655) );
  NAND2XL U1640 ( .A(n2656), .B(n2661), .Y(n2663) );
  NAND2XL U1641 ( .A(n144), .B(n2649), .Y(n2653) );
  NAND2XL U1642 ( .A(n2645), .B(n2644), .Y(n2649) );
  NOR2XL U1643 ( .A(n2646), .B(n2642), .Y(n2643) );
  INVXL U1644 ( .A(n2654), .Y(n2646) );
  INVXL U1645 ( .A(n2642), .Y(n2648) );
  NAND2BXL U1646 ( .AN(n2635), .B(n2638), .Y(n2644) );
  NAND2XL U1647 ( .A(n2631), .B(n2633), .Y(n2638) );
  NAND2XL U1648 ( .A(n145), .B(n2629), .Y(n2633) );
  NAND2XL U1649 ( .A(n2627), .B(n2632), .Y(n2626) );
  NOR2XL U1650 ( .A(n2628), .B(n2627), .Y(n2625) );
  NAND2BXL U1651 ( .AN(n2616), .B(n2621), .Y(n2618) );
  NAND2XL U1652 ( .A(n2615), .B(n2614), .Y(n2621) );
  NAND2XL U1653 ( .A(n2611), .B(n2610), .Y(n2614) );
  NAND2XL U1654 ( .A(n2608), .B(n2612), .Y(n2607) );
  NOR2XL U1655 ( .A(n2609), .B(n2608), .Y(n2606) );
  INVXL U1656 ( .A(n2613), .Y(n2609) );
  NAND2BXL U1657 ( .AN(n2597), .B(n2602), .Y(n2599) );
  NAND2XL U1658 ( .A(n2596), .B(n2595), .Y(n2602) );
  NAND2XL U1659 ( .A(n143), .B(n2591), .Y(n2595) );
  NAND2XL U1660 ( .A(n2589), .B(n2593), .Y(n2588) );
  NOR2XL U1661 ( .A(n2590), .B(n2589), .Y(n2587) );
  NAND2BXL U1662 ( .AN(n2578), .B(n2583), .Y(n2580) );
  NAND2XL U1663 ( .A(n2577), .B(n2576), .Y(n2583) );
  NAND2XL U1664 ( .A(n2573), .B(n2572), .Y(n2576) );
  NAND2XL U1665 ( .A(n2570), .B(n2574), .Y(n2569) );
  NOR2XL U1666 ( .A(n2571), .B(n2570), .Y(n2568) );
  NAND2BXL U1667 ( .AN(n149), .B(n2564), .Y(n2561) );
  NAND2XL U1668 ( .A(n2558), .B(n2557), .Y(n2564) );
  NAND2XL U1669 ( .A(n2554), .B(n2553), .Y(n2557) );
  NAND2XL U1670 ( .A(n2551), .B(n2555), .Y(n2550) );
  NOR2XL U1671 ( .A(n2552), .B(n2551), .Y(n2549) );
  NAND2XL U1672 ( .A(n2543), .B(n2544), .Y(n2553) );
  NAND2BXL U1673 ( .AN(n2542), .B(n2546), .Y(n2544) );
  NAND2XL U1674 ( .A(n2541), .B(n2540), .Y(n2546) );
  NAND2XL U1675 ( .A(n2537), .B(n2536), .Y(n2540) );
  NAND2XL U1676 ( .A(n2534), .B(n2538), .Y(n2533) );
  NOR2XL U1677 ( .A(n2535), .B(n2534), .Y(n2532) );
  NAND2BXL U1678 ( .AN(n2523), .B(n2528), .Y(n2525) );
  NOR2XL U1679 ( .A(n2519), .B(n2515), .Y(n2517) );
  AOI211XL U1680 ( .A0(n2514), .A1(n2860), .B0(n2867), .C0(n2513), .Y(n2677)
         );
  NOR2XL U1681 ( .A(n2512), .B(n2514), .Y(n2513) );
  XOR2XL U1682 ( .A(n2509), .B(n2508), .Y(n2510) );
  NAND3XL U1683 ( .A(n2506), .B(N1826), .C(n232), .Y(n2504) );
  NAND3XL U1684 ( .A(n2498), .B(n2500), .C(n2503), .Y(n2499) );
  AND2XL U1685 ( .A(n2497), .B(n2496), .Y(n2498) );
  NAND2XL U1686 ( .A(n2500), .B(n2503), .Y(n2492) );
  NOR2XL U1687 ( .A(n2495), .B(n2494), .Y(n2491) );
  NOR2XL U1688 ( .A(n2486), .B(n164), .Y(n2487) );
  INVXL U1689 ( .A(n2495), .Y(n2484) );
  INVXL U1690 ( .A(n2479), .Y(n2475) );
  NAND3XL U1691 ( .A(n2480), .B(n2474), .C(n2481), .Y(n2479) );
  INVXL U1692 ( .A(n2481), .Y(n2470) );
  INVXL U1693 ( .A(n2480), .Y(n2471) );
  INVXL U1694 ( .A(n2465), .Y(n2459) );
  NOR2XL U1695 ( .A(work_cntr[4]), .B(n2477), .Y(n2460) );
  NAND3XL U1696 ( .A(n2466), .B(n2458), .C(n2461), .Y(n2474) );
  NAND3XL U1697 ( .A(n2463), .B(n2462), .C(n2457), .Y(n2461) );
  INVXL U1698 ( .A(n2455), .Y(n2462) );
  INVXL U1699 ( .A(n2458), .Y(n2468) );
  NOR2XL U1700 ( .A(work_cntr[7]), .B(n2464), .Y(n2448) );
  NAND3XL U1701 ( .A(n2452), .B(n2453), .C(n2449), .Y(n2457) );
  NAND2XL U1702 ( .A(n2451), .B(n2441), .Y(n2445) );
  NAND3XL U1703 ( .A(n2437), .B(n2431), .C(n2434), .Y(n2441) );
  NAND3XL U1704 ( .A(n2436), .B(n2430), .C(n2435), .Y(n2434) );
  INVXL U1705 ( .A(n2431), .Y(n2439) );
  INVXL U1706 ( .A(n2435), .Y(n2428) );
  NAND2XL U1707 ( .A(n2476), .B(n2414), .Y(n2416) );
  NAND2XL U1708 ( .A(n2422), .B(n2412), .Y(n2430) );
  AOI32XL U1709 ( .A0(n2404), .A1(n2403), .A2(n2402), .B0(n2401), .B1(n2403), 
        .Y(n2407) );
  NAND2BXL U1710 ( .AN(n2400), .B(n2401), .Y(n2403) );
  INVXL U1711 ( .A(n2425), .Y(n2412) );
  NOR2XL U1712 ( .A(n2418), .B(n2409), .Y(n2410) );
  INVXL U1713 ( .A(n2396), .Y(n2401) );
  NOR2XL U1714 ( .A(work_cntr[15]), .B(n2393), .Y(n2395) );
  NAND2XL U1715 ( .A(n2391), .B(n2390), .Y(n2404) );
  NAND2BXL U1716 ( .AN(n2402), .B(n2392), .Y(n2398) );
  NAND2XL U1717 ( .A(n2385), .B(work_cntr[19]), .Y(n2384) );
  NAND2XL U1718 ( .A(n2383), .B(n2432), .Y(n2394) );
  INVXL U1719 ( .A(n2433), .Y(n2432) );
  INVXL U1720 ( .A(n2399), .Y(n2406) );
  NOR2XL U1721 ( .A(n2374), .B(n2373), .Y(n2375) );
  AOI211XL U1722 ( .A0(n2372), .A1(n2371), .B0(n2370), .C0(n2369), .Y(n2373)
         );
  NOR2XL U1723 ( .A(n2372), .B(n2371), .Y(n2369) );
  NAND2XL U1724 ( .A(n2368), .B(n2367), .Y(n2370) );
  AOI211XL U1725 ( .A0(n2362), .A1(n2361), .B0(n2360), .C0(n2359), .Y(n2368)
         );
  NOR2XL U1726 ( .A(n2358), .B(n2362), .Y(n2359) );
  NOR2XL U1727 ( .A(n2353), .B(n2352), .Y(n2374) );
  NOR2XL U1728 ( .A(n2351), .B(n2350), .Y(n2376) );
  NAND2XL U1729 ( .A(n2353), .B(n2352), .Y(n2377) );
  NAND2XL U1730 ( .A(n2351), .B(n2350), .Y(n2352) );
  INVXL U1731 ( .A(n2362), .Y(n2348) );
  INVXL U1732 ( .A(n2337), .Y(n2339) );
  NOR4BXL U1733 ( .AN(n2361), .B(n2341), .C(n2357), .D(n2363), .Y(n2349) );
  NOR2XL U1734 ( .A(n2331), .B(n2330), .Y(n2332) );
  INVXL U1735 ( .A(n2351), .Y(next_work_cntr[0]) );
  INVXL U1736 ( .A(n2327), .Y(n2340) );
  NAND2XL U1737 ( .A(n2347), .B(n2346), .Y(n2326) );
  NAND2XL U1738 ( .A(n2343), .B(n2320), .Y(n2321) );
  INVXL U1739 ( .A(n2338), .Y(n2320) );
  NAND2XL U1740 ( .A(n2317), .B(n2316), .Y(n2338) );
  NAND2XL U1741 ( .A(n2371), .B(n2354), .Y(n2329) );
  INVXL U1742 ( .A(n2299), .Y(n2325) );
  NOR4XL U1743 ( .A(next_work_cntr[2]), .B(n2292), .C(n2291), .D(n2331), .Y(
        n2293) );
  INVXL U1744 ( .A(n2307), .Y(n2292) );
  INVXL U1745 ( .A(n2343), .Y(n2301) );
  INVXL U1746 ( .A(n2334), .Y(n2366) );
  INVXL U1747 ( .A(n2283), .Y(n2286) );
  NAND2XL U1748 ( .A(n2280), .B(n2287), .Y(n2281) );
  NAND2XL U1749 ( .A(n2279), .B(n2285), .Y(n2287) );
  NAND2XL U1750 ( .A(n2307), .B(n2306), .Y(n2310) );
  INVXL U1751 ( .A(n2271), .Y(n2274) );
  NAND2BXL U1752 ( .AN(n2298), .B(n211), .Y(n2268) );
  NAND4BXL U1753 ( .AN(n2288), .B(n2279), .C(n2307), .D(n2282), .Y(n2275) );
  NAND2XL U1754 ( .A(n2265), .B(n2264), .Y(n2283) );
  INVXL U1755 ( .A(n2256), .Y(n2257) );
  INVXL U1756 ( .A(n2250), .Y(n2253) );
  NOR2XL U1757 ( .A(n2245), .B(n2244), .Y(n2247) );
  NAND4BXL U1758 ( .AN(n2255), .B(n2254), .C(n2266), .D(n2269), .Y(n2249) );
  NAND2BXL U1759 ( .AN(n2234), .B(n2233), .Y(n2235) );
  NAND2XL U1760 ( .A(n2256), .B(n2259), .Y(n2233) );
  INVXL U1761 ( .A(n2265), .Y(next_work_cntr[4]) );
  NAND2XL U1762 ( .A(n2259), .B(n2282), .Y(n2255) );
  NAND2XL U1763 ( .A(n2251), .B(n2250), .Y(n2223) );
  NAND2XL U1764 ( .A(n2252), .B(n2246), .Y(n2251) );
  NAND2XL U1765 ( .A(n2222), .B(n2225), .Y(n2232) );
  NAND2XL U1766 ( .A(n2207), .B(n2206), .Y(n2208) );
  INVXL U1767 ( .A(n2634), .Y(n2628) );
  AND2XL U1768 ( .A(n2204), .B(next_work_cntr[6]), .Y(n2221) );
  INVXL U1769 ( .A(n2199), .Y(n2197) );
  AOI21XL U1770 ( .A0(n2191), .A1(n2190), .B0(n2189), .Y(n2192) );
  NAND4BXL U1771 ( .AN(n2215), .B(n2212), .C(n2205), .D(n2188), .Y(n2195) );
  NAND2BXL U1772 ( .AN(n2236), .B(n166), .Y(n2217) );
  INVXL U1773 ( .A(n2186), .Y(n2228) );
  AOI211XL U1774 ( .A0(n2185), .A1(n2184), .B0(n2183), .C0(n2182), .Y(n2186)
         );
  NOR2XL U1775 ( .A(n2185), .B(n2184), .Y(n2182) );
  INVXL U1776 ( .A(n2181), .Y(n2184) );
  NAND2XL U1777 ( .A(n2203), .B(n2222), .Y(n2227) );
  AND2XL U1778 ( .A(n166), .B(n2229), .Y(n2175) );
  INVXL U1779 ( .A(n2187), .Y(n2229) );
  NAND2XL U1780 ( .A(n2181), .B(n2183), .Y(n2187) );
  OAI2BB2XL U1781 ( .B0(n2169), .B1(n2168), .A0N(n2169), .A1N(n2168), .Y(n2231) );
  NOR2XL U1782 ( .A(n136), .B(n2165), .Y(n2167) );
  INVXL U1783 ( .A(n2164), .Y(n2173) );
  INVXL U1784 ( .A(n2160), .Y(n2163) );
  INVXL U1785 ( .A(n2152), .Y(n2158) );
  NAND3XL U1786 ( .A(n2172), .B(n2203), .C(n2177), .Y(n2150) );
  AOI211XL U1787 ( .A0(next_work_cntr[12]), .A1(n2147), .B0(n2146), .C0(n2149), 
        .Y(n2148) );
  NAND2XL U1788 ( .A(n2145), .B(n2144), .Y(n2147) );
  INVXL U1789 ( .A(n2153), .Y(next_work_cntr[12]) );
  NAND2XL U1790 ( .A(n2169), .B(n2166), .Y(n2164) );
  NAND2XL U1791 ( .A(n2161), .B(n2160), .Y(n2136) );
  NAND2XL U1792 ( .A(n2141), .B(n2162), .Y(n2161) );
  NOR2XL U1793 ( .A(n2140), .B(n2139), .Y(n2130) );
  NOR2XL U1794 ( .A(next_work_cntr[16]), .B(n2127), .Y(n2131) );
  NAND2XL U1795 ( .A(n2155), .B(n2149), .Y(n2152) );
  INVXL U1796 ( .A(n2123), .Y(n2144) );
  NAND2XL U1797 ( .A(n2169), .B(n2181), .Y(n2151) );
  NAND2XL U1798 ( .A(n2169), .B(n2120), .Y(n2121) );
  NAND2XL U1799 ( .A(n2146), .B(n2116), .Y(n2117) );
  NAND2XL U1800 ( .A(n2114), .B(next_work_cntr[19]), .Y(n2135) );
  INVXL U1801 ( .A(next_work_cntr[16]), .Y(n2113) );
  AOI32XL U1802 ( .A0(n2111), .A1(n318), .A2(n2790), .B0(si_sel), .B1(n2110), 
        .Y(n2680) );
  AOI211XL U1803 ( .A0(n2109), .A1(n2108), .B0(n2351), .C0(n2107), .Y(n2110)
         );
  NOR2XL U1804 ( .A(n2106), .B(n2109), .Y(n2107) );
  NOR2XL U1805 ( .A(n2105), .B(n2104), .Y(n2106) );
  INVXL U1806 ( .A(n2091), .Y(n2092) );
  INVXL U1807 ( .A(n2100), .Y(n2093) );
  INVXL U1808 ( .A(n2090), .Y(n2096) );
  NOR3XL U1809 ( .A(N1826), .B(n2089), .C(n317), .Y(n2097) );
  NOR2XL U1810 ( .A(n2079), .B(n2078), .Y(n2081) );
  OAI211XL U1811 ( .A0(n2089), .A1(n2085), .B0(n2090), .C0(n2087), .Y(n2082)
         );
  NAND2XL U1812 ( .A(n2077), .B(n2076), .Y(n2087) );
  NAND2XL U1813 ( .A(n263), .B(n316), .Y(n2085) );
  XNOR2XL U1814 ( .A(n2072), .B(n2070), .Y(n2073) );
  INVXL U1815 ( .A(n2083), .Y(n2069) );
  NAND2XL U1816 ( .A(n2063), .B(n2062), .Y(n2064) );
  NAND2BXL U1817 ( .AN(n2072), .B(n2070), .Y(n2062) );
  NOR2XL U1818 ( .A(n2071), .B(n2072), .Y(n2066) );
  NOR2XL U1819 ( .A(n2053), .B(n2058), .Y(n2056) );
  NAND2XL U1820 ( .A(n2065), .B(n2054), .Y(n2053) );
  INVXL U1821 ( .A(n2046), .Y(n2047) );
  NAND2BXL U1822 ( .AN(n2057), .B(n2045), .Y(n2051) );
  NOR3XL U1823 ( .A(n2044), .B(n2043), .C(n2057), .Y(n2052) );
  INVXL U1824 ( .A(n2041), .Y(n2042) );
  INVXL U1825 ( .A(n2049), .Y(n2043) );
  AND2XL U1826 ( .A(n2035), .B(n2034), .Y(n2048) );
  NAND3XL U1827 ( .A(n2035), .B(n2049), .C(n2030), .Y(n2037) );
  AOI211XL U1828 ( .A0(n2028), .A1(n2032), .B0(n2022), .C0(n2026), .Y(n2023)
         );
  INVXL U1829 ( .A(n2019), .Y(n2022) );
  OAI211XL U1830 ( .A0(n2013), .A1(n2021), .B0(n2012), .C0(n2019), .Y(n2014)
         );
  INVXL U1831 ( .A(n2017), .Y(n2015) );
  NAND2XL U1832 ( .A(n2012), .B(n2013), .Y(n2017) );
  XOR2XL U1833 ( .A(n168), .B(n2010), .Y(n2016) );
  NOR2XL U1834 ( .A(n168), .B(n1999), .Y(n2006) );
  INVXL U1835 ( .A(n1999), .Y(n2010) );
  NAND2XL U1836 ( .A(n1997), .B(n1996), .Y(n1999) );
  NAND2XL U1837 ( .A(n1989), .B(n2001), .Y(n1995) );
  NAND3XL U1838 ( .A(n1989), .B(n167), .C(n1997), .Y(n2004) );
  OAI2BB2XL U1839 ( .B0(n1988), .B1(n1987), .A0N(n1988), .A1N(n1987), .Y(n2011) );
  INVXL U1840 ( .A(n169), .Y(n1989) );
  AND2XL U1841 ( .A(n1991), .B(n1983), .Y(n1980) );
  NAND4XL U1842 ( .A(n1972), .B(n1971), .C(n1970), .D(n1974), .Y(n1973) );
  NAND2XL U1843 ( .A(n1979), .B(n1978), .Y(n1991) );
  XOR2XL U1844 ( .A(n1967), .B(n1974), .Y(n1968) );
  NAND2XL U1845 ( .A(n1972), .B(n1961), .Y(n1962) );
  INVXL U1846 ( .A(n1963), .Y(n1961) );
  NAND4XL U1847 ( .A(n1955), .B(n2521), .C(n2520), .D(n2522), .Y(n2108) );
  NOR4XL U1848 ( .A(n2571), .B(n2112), .C(n1954), .D(n2527), .Y(n1955) );
  INVXL U1849 ( .A(n2526), .Y(n2527) );
  NAND4XL U1850 ( .A(n1953), .B(n2594), .C(n2562), .D(n2539), .Y(n1954) );
  INVXL U1851 ( .A(n2535), .Y(n2539) );
  AOI211XL U1852 ( .A0(n1952), .A1(n1951), .B0(n1950), .C0(n1949), .Y(n1953)
         );
  NAND4XL U1853 ( .A(n2600), .B(n2613), .C(n2619), .D(n2634), .Y(n1949) );
  INVXL U1854 ( .A(n2562), .Y(n2563) );
  NAND2XL U1855 ( .A(n1000), .B(work_cntr[12]), .Y(n999) );
  INVXL U1856 ( .A(n1001), .Y(n1000) );
  NAND2XL U1857 ( .A(write_addr[16]), .B(n134), .Y(n372) );
  NAND2XL U1858 ( .A(n134), .B(\next_write_addr_w[0] ), .Y(n377) );
  NAND2XL U1859 ( .A(n134), .B(write_addr[5]), .Y(n361) );
  NAND2XL U1860 ( .A(n135), .B(n713), .Y(n357) );
  NAND2XL U1861 ( .A(n134), .B(write_addr[6]), .Y(n362) );
  NAND2XL U1862 ( .A(write_addr[8]), .B(n134), .Y(n374) );
  INVXL U1863 ( .A(n2830), .Y(n373) );
  INVXL U1864 ( .A(n582), .Y(n375) );
  MXI2XL U1865 ( .A(n703), .B(n288), .S0(n134), .Y(n481) );
  MXI2XL U1866 ( .A(n2850), .B(n292), .S0(n134), .Y(n443) );
  NAND2XL U1867 ( .A(n134), .B(write_addr[3]), .Y(n359) );
  NAND2XL U1868 ( .A(n134), .B(write_addr[7]), .Y(n363) );
  NOR4XL U1869 ( .A(n2859), .B(n1793), .C(n2684), .D(n318), .Y(n1794) );
  NOR4XL U1870 ( .A(N196), .B(n1792), .C(n1791), .D(n1790), .Y(n1793) );
  OAI211XL U1871 ( .A0(n2378), .A1(n1777), .B0(n1779), .C0(n2497), .Y(n1764)
         );
  NOR2XL U1872 ( .A(n1763), .B(n1765), .Y(n1766) );
  AOI211XL U1873 ( .A0(n1759), .A1(n1758), .B0(n1767), .C0(n1757), .Y(n1760)
         );
  NOR2XL U1874 ( .A(n1759), .B(n1758), .Y(n1757) );
  NAND2XL U1875 ( .A(n1748), .B(n1747), .Y(n1752) );
  INVXL U1876 ( .A(n1765), .Y(n1755) );
  INVXL U1877 ( .A(n1741), .Y(n1748) );
  INVXL U1878 ( .A(n1747), .Y(n1744) );
  NAND2XL U1879 ( .A(n1726), .B(n1725), .Y(n1729) );
  INVXL U1880 ( .A(n1724), .Y(n1732) );
  OAI211XL U1881 ( .A0(n137), .A1(n1717), .B0(n1719), .C0(n1720), .Y(n1718) );
  INVXL U1882 ( .A(n1716), .Y(n1717) );
  AND2XL U1883 ( .A(n153), .B(n1710), .Y(n1700) );
  NOR2BXL U1884 ( .AN(n1706), .B(n1698), .Y(n1711) );
  NOR2XL U1885 ( .A(n1698), .B(n1699), .Y(n1703) );
  INVXL U1886 ( .A(n1707), .Y(n1698) );
  INVXL U1887 ( .A(n1688), .Y(n1691) );
  INVXL U1888 ( .A(n1684), .Y(n1683) );
  INVXL U1889 ( .A(n1677), .Y(n1679) );
  NAND2XL U1890 ( .A(n1676), .B(n1675), .Y(n1681) );
  AOI211XL U1891 ( .A0(n1685), .A1(n1686), .B0(n1674), .C0(n1673), .Y(n1682)
         );
  NOR2XL U1892 ( .A(work_cntr[12]), .B(n1689), .Y(n1672) );
  NOR2BXL U1893 ( .AN(n1686), .B(n1673), .Y(n1693) );
  INVXL U1894 ( .A(n1663), .Y(n1666) );
  NAND2XL U1895 ( .A(n1687), .B(n1669), .Y(n1677) );
  NAND2XL U1896 ( .A(n1661), .B(n1660), .Y(n1675) );
  NOR2XL U1897 ( .A(n1657), .B(n1656), .Y(n1658) );
  NAND4XL U1898 ( .A(n1651), .B(n1650), .C(n1665), .D(n1653), .Y(n1652) );
  NOR2XL U1899 ( .A(n1651), .B(n1656), .Y(n1648) );
  INVXL U1900 ( .A(n1647), .Y(n1656) );
  NOR2XL U1901 ( .A(work_cntr[15]), .B(n1655), .Y(n1646) );
  INVXL U1902 ( .A(n1651), .Y(n1657) );
  AOI222XL U1903 ( .A0(n729), .A1(\C159/DATA3_19 ), .B0(n746), .B1(
        global_cntr[19]), .C0(n311), .C1(N1366), .Y(\im_a[19]_BAR ) );
  INVXL U1904 ( .A(n1785), .Y(n726) );
  NOR2XL U1905 ( .A(n1786), .B(\sftr_n[0]_BAR ), .Y(n727) );
  NOR2BXL U1906 ( .AN(curr_photo_addr[19]), .B(n313), .Y(\C1/Z_19 ) );
  OAI211XL U1907 ( .A0(n710), .A1(n158), .B0(n571), .C0(n570), .Y(n572) );
  AOI211XL U1908 ( .A0(n723), .A1(n713), .B0(n712), .C0(n711), .Y(n714) );
  OAI211XL U1909 ( .A0(n716), .A1(n710), .B0(n709), .C0(n708), .Y(n711) );
  NAND2XL U1910 ( .A(n707), .B(write_addr[2]), .Y(n708) );
  AOI211XL U1911 ( .A0(n720), .A1(write_addr[2]), .B0(n706), .C0(n705), .Y(
        n709) );
  NOR2XL U1912 ( .A(n2834), .B(n717), .Y(n706) );
  NOR2XL U1913 ( .A(n703), .B(n715), .Y(n712) );
  AOI211XL U1914 ( .A0(write_addr[8]), .A1(n2855), .B0(n2783), .C0(n1824), .Y(
        n376) );
  AOI32XL U1915 ( .A0(n1823), .A1(n1822), .A2(write_addr[8]), .B0(n2707), .B1(
        n1894), .Y(n1824) );
  INVXL U1916 ( .A(n1894), .Y(n1822) );
  OAI211XL U1917 ( .A0(n701), .A1(n700), .B0(n699), .C0(n698), .Y(n702) );
  NAND2XL U1918 ( .A(n697), .B(n713), .Y(n698) );
  AOI211XL U1919 ( .A0(n696), .A1(n722), .B0(n695), .C0(n694), .Y(n699) );
  AOI21XL U1920 ( .A0(n720), .A1(write_addr[3]), .B0(n692), .Y(n693) );
  NOR2XL U1921 ( .A(n721), .B(n289), .Y(n695) );
  NAND2XL U1922 ( .A(n1931), .B(n288), .Y(n358) );
  OAI211XL U1923 ( .A0(n1929), .A1(n1903), .B0(n310), .C0(n1902), .Y(n1904) );
  NAND2XL U1924 ( .A(n1929), .B(n1903), .Y(n1902) );
  INVXL U1925 ( .A(n1911), .Y(n1901) );
  AOI211XL U1926 ( .A0(n723), .A1(n690), .B0(n689), .C0(n688), .Y(n691) );
  OAI211XL U1927 ( .A0(n741), .A1(n721), .B0(n687), .C0(n686), .Y(n688) );
  NAND2XL U1928 ( .A(n696), .B(n713), .Y(n686) );
  AOI211XL U1929 ( .A0(n720), .A1(write_addr[4]), .B0(n685), .C0(n684), .Y(
        n687) );
  NOR2XL U1930 ( .A(n717), .B(n683), .Y(n685) );
  INVXL U1931 ( .A(n707), .Y(n721) );
  NOR2XL U1932 ( .A(n701), .B(n715), .Y(n689) );
  AOI211XL U1933 ( .A0(n697), .A1(n690), .B0(n681), .C0(n680), .Y(n682) );
  OAI211XL U1934 ( .A0(n701), .A1(n710), .B0(n679), .C0(n678), .Y(n680) );
  NAND2XL U1935 ( .A(n707), .B(write_addr[5]), .Y(n678) );
  AOI211XL U1936 ( .A0(n720), .A1(write_addr[5]), .B0(n677), .C0(n676), .Y(
        n679) );
  NOR2XL U1937 ( .A(n717), .B(n2838), .Y(n677) );
  NOR2XL U1938 ( .A(n675), .B(n700), .Y(n681) );
  NOR2BXL U1939 ( .AN(curr_photo_addr[5]), .B(n313), .Y(n734) );
  AOI211XL U1940 ( .A0(n696), .A1(n690), .B0(n672), .C0(n671), .Y(n673) );
  OAI211XL U1941 ( .A0(n2839), .A1(n717), .B0(n670), .C0(n669), .Y(n671) );
  NAND2XL U1942 ( .A(n707), .B(write_addr[6]), .Y(n669) );
  AOI21XL U1943 ( .A0(n720), .A1(write_addr[6]), .B0(n668), .Y(n670) );
  NOR2XL U1944 ( .A(n675), .B(n715), .Y(n672) );
  NOR2BXL U1945 ( .AN(curr_photo_addr[6]), .B(n313), .Y(n735) );
  AOI211XL U1946 ( .A0(n723), .A1(n666), .B0(n665), .C0(n664), .Y(n667) );
  OAI211XL U1947 ( .A0(n675), .A1(n710), .B0(n663), .C0(n662), .Y(n664) );
  NAND2XL U1948 ( .A(n707), .B(write_addr[7]), .Y(n662) );
  AOI211XL U1949 ( .A0(n720), .A1(write_addr[7]), .B0(n661), .C0(n660), .Y(
        n663) );
  NOR2XL U1950 ( .A(n2840), .B(n717), .Y(n661) );
  NOR2XL U1951 ( .A(n2845), .B(n715), .Y(n665) );
  AOI211XL U1952 ( .A0(n697), .A1(n666), .B0(n658), .C0(n657), .Y(n659) );
  AOI211XL U1953 ( .A0(\C158/DATA2_7 ), .A1(n720), .B0(n655), .C0(n654), .Y(
        n656) );
  AOI21XL U1954 ( .A0(n2843), .A1(n2842), .B0(n2841), .Y(n2844) );
  NOR2XL U1955 ( .A(write_addr[9]), .B(n651), .Y(n655) );
  XOR2XL U1956 ( .A(\C1/Z_7 ), .B(write_addr[9]), .Y(\C158/DATA2_7 ) );
  NOR2XL U1957 ( .A(n650), .B(n700), .Y(n658) );
  INVXL U1958 ( .A(n2852), .Y(n666) );
  NOR2BXL U1959 ( .AN(curr_photo_addr[8]), .B(n313), .Y(\C1/Z_8 ) );
  AOI211XL U1960 ( .A0(n723), .A1(n648), .B0(n647), .C0(n646), .Y(n649) );
  OAI211XL U1961 ( .A0(n2852), .A1(n710), .B0(n645), .C0(n644), .Y(n646) );
  NAND2XL U1962 ( .A(n720), .B(\C158/DATA2_8 ), .Y(n644) );
  AOI211XL U1963 ( .A0(n707), .A1(write_addr[10]), .B0(n643), .C0(n642), .Y(
        n645) );
  AOI211XL U1964 ( .A0(n2849), .A1(n292), .B0(n717), .C0(n2848), .Y(n643) );
  NAND2XL U1965 ( .A(n2847), .B(write_addr[9]), .Y(n2849) );
  NAND2XL U1966 ( .A(n744), .B(n1825), .Y(n1944) );
  NOR2XL U1967 ( .A(n2846), .B(n715), .Y(n647) );
  NOR2BXL U1968 ( .AN(curr_photo_addr[9]), .B(n313), .Y(\C1/Z_9 ) );
  NOR2BXL U1969 ( .AN(curr_photo_addr[10]), .B(n313), .Y(\C1/Z_10 ) );
  AOI211XL U1970 ( .A0(n697), .A1(n648), .B0(n640), .C0(n639), .Y(n641) );
  OAI211XL U1971 ( .A0(n2846), .A1(n710), .B0(n638), .C0(n637), .Y(n639) );
  NAND2XL U1972 ( .A(n720), .B(\C158/DATA2_10 ), .Y(n637) );
  AOI211XL U1973 ( .A0(n636), .A1(write_addr[8]), .B0(n635), .C0(n634), .Y(
        n638) );
  NAND2XL U1974 ( .A(n652), .B(write_addr[10]), .Y(n633) );
  NOR4XL U1975 ( .A(n717), .B(write_addr[12]), .C(n2816), .D(n223), .Y(n635)
         );
  NOR2XL U1976 ( .A(n632), .B(n700), .Y(n640) );
  INVXL U1977 ( .A(n2850), .Y(n648) );
  AOI211XL U1978 ( .A0(n2858), .A1(n697), .B0(n630), .C0(n629), .Y(n631) );
  AOI211XL U1979 ( .A0(\C158/DATA2_11 ), .A1(n720), .B0(n627), .C0(n626), .Y(
        n628) );
  AOI211XL U1980 ( .A0(n2823), .A1(n296), .B0(n625), .C0(\sftr_n[0]_BAR ), .Y(
        n627) );
  AND3XL U1981 ( .A(write_addr[13]), .B(n2819), .C(n2818), .Y(n625) );
  NAND2XL U1982 ( .A(n2826), .B(n297), .Y(n2818) );
  INVXL U1983 ( .A(n2856), .Y(n2819) );
  NOR2XL U1984 ( .A(n223), .B(n2816), .Y(n2817) );
  INVXL U1985 ( .A(n2848), .Y(n2816) );
  NOR2XL U1986 ( .A(n624), .B(n700), .Y(n630) );
  NOR2BXL U1987 ( .AN(curr_photo_addr[12]), .B(n313), .Y(\C1/Z_12 ) );
  AOI211XL U1988 ( .A0(n720), .A1(\C158/DATA2_12 ), .B0(n621), .C0(n620), .Y(
        n622) );
  OAI211XL U1989 ( .A0(n619), .A1(n700), .B0(n618), .C0(n617), .Y(n620) );
  NAND3XL U1990 ( .A(n616), .B(n2821), .C(n740), .Y(n617) );
  NOR2XL U1991 ( .A(n2850), .B(n710), .Y(n621) );
  AOI211XL U1992 ( .A0(n292), .A1(n2714), .B0(n2713), .C0(n2783), .Y(n2716) );
  OAI211XL U1993 ( .A0(n624), .A1(n715), .B0(n614), .C0(n613), .Y(n615) );
  NAND2XL U1994 ( .A(n696), .B(n2858), .Y(n613) );
  AOI211XL U1995 ( .A0(n2756), .A1(n2755), .B0(n2762), .C0(n2783), .Y(n2757)
         );
  XOR2XL U1996 ( .A(\intadd_3/B[8] ), .B(\intadd_3/n3 ), .Y(\intadd_3/SUM[8] )
         );
  AOI211XL U1997 ( .A0(\C158/DATA2_13 ), .A1(n720), .B0(n612), .C0(n611), .Y(
        n614) );
  OAI211XL U1998 ( .A0(n223), .A1(n704), .B0(n610), .C0(n609), .Y(n611) );
  OAI211XL U1999 ( .A0(n2821), .A1(n299), .B0(n740), .C0(n608), .Y(n609) );
  NAND2XL U2000 ( .A(write_addr[13]), .B(n652), .Y(n610) );
  NOR2XL U2001 ( .A(n700), .B(n607), .Y(n612) );
  AOI211XL U2002 ( .A0(n720), .A1(\C158/DATA2_14 ), .B0(n605), .C0(n604), .Y(
        n606) );
  OAI211XL U2003 ( .A0(n603), .A1(n700), .B0(n602), .C0(n601), .Y(n604) );
  OAI211XL U2004 ( .A0(write_addr[16]), .A1(n600), .B0(n2825), .C0(n740), .Y(
        n601) );
  NOR2XL U2005 ( .A(n2823), .B(n2824), .Y(n600) );
  NOR2XL U2006 ( .A(n632), .B(n710), .Y(n605) );
  OAI211XL U2007 ( .A0(n624), .A1(n710), .B0(n597), .C0(n596), .Y(n598) );
  NAND2XL U2008 ( .A(n720), .B(\C158/DATA2_15 ), .Y(n596) );
  AOI211XL U2009 ( .A0(n159), .A1(n723), .B0(n595), .C0(n594), .Y(n597) );
  OAI211XL U2010 ( .A0(n607), .A1(n715), .B0(n593), .C0(n592), .Y(n594) );
  OAI211XL U2011 ( .A0(n2825), .A1(n283), .B0(n740), .C0(n591), .Y(n592) );
  INVXL U2012 ( .A(n2853), .Y(n2826) );
  NAND2XL U2013 ( .A(n652), .B(write_addr[15]), .Y(n593) );
  NOR2XL U2014 ( .A(n704), .B(n296), .Y(n595) );
  INVXL U2015 ( .A(n2828), .Y(n624) );
  AOI211XL U2016 ( .A0(n2766), .A1(n2765), .B0(n2773), .C0(n2783), .Y(n2767)
         );
  AND2XL U2017 ( .A(\intadd_3/A[9] ), .B(n245), .Y(n246) );
  NAND2XL U2018 ( .A(n1911), .B(n1910), .Y(n1912) );
  NOR2XL U2019 ( .A(n1911), .B(n1910), .Y(n1913) );
  INVXL U2020 ( .A(n1908), .Y(n1898) );
  NAND2XL U2021 ( .A(n1897), .B(n174), .Y(n1899) );
  INVXL U2022 ( .A(n1892), .Y(n1897) );
  AOI21XL U2023 ( .A0(n1937), .A1(n1922), .B0(n1935), .Y(\intadd_3/B[0] ) );
  INVXL U2024 ( .A(n1918), .Y(\intadd_3/A[0] ) );
  INVXL U2025 ( .A(n1930), .Y(\intadd_3/B[1] ) );
  NAND2XL U2026 ( .A(n1909), .B(n1936), .Y(n1927) );
  NAND2BXL U2027 ( .AN(n1887), .B(n1886), .Y(n1888) );
  AOI211XL U2028 ( .A0(n1929), .A1(n1880), .B0(n1879), .C0(n1878), .Y(n1881)
         );
  NOR2XL U2029 ( .A(n1929), .B(n1880), .Y(n1874) );
  NAND2BXL U2030 ( .AN(n1868), .B(n1887), .Y(n1884) );
  AND2XL U2031 ( .A(n1905), .B(n174), .Y(n1920) );
  INVXL U2032 ( .A(n1869), .Y(n1872) );
  INVXL U2033 ( .A(n1867), .Y(n1863) );
  NAND2XL U2034 ( .A(n1861), .B(n1936), .Y(n1867) );
  INVXL U2035 ( .A(n1875), .Y(n1860) );
  INVXL U2036 ( .A(n1851), .Y(n1854) );
  NAND2XL U2037 ( .A(n1871), .B(n1862), .Y(n1870) );
  NAND2XL U2038 ( .A(n1864), .B(n1861), .Y(n1862) );
  AND3XL U2039 ( .A(n1845), .B(n1843), .C(n1941), .Y(n1841) );
  INVXL U2040 ( .A(n1836), .Y(n1839) );
  NAND2XL U2041 ( .A(n1853), .B(n1840), .Y(n1852) );
  NAND3XL U2042 ( .A(n1845), .B(n1842), .C(n1843), .Y(n1840) );
  NAND2XL U2043 ( .A(n1850), .B(n1847), .Y(n1843) );
  AND3XL U2044 ( .A(n1833), .B(n1834), .C(n2704), .Y(n1827) );
  INVXL U2045 ( .A(n1019), .Y(n1022) );
  NAND2XL U2046 ( .A(n1838), .B(n1826), .Y(n1837) );
  NAND3XL U2047 ( .A(n1828), .B(n1833), .C(n1834), .Y(n1826) );
  AND3XL U2048 ( .A(n1014), .B(n1012), .C(next_cr_x[5]), .Y(n1010) );
  XOR2XL U2049 ( .A(n307), .B(next_cr_x[6]), .Y(\DP_OP_589J1_125_1438/n26 ) );
  XOR2XL U2050 ( .A(n174), .B(next_cr_x[5]), .Y(n307) );
  MXI2XL U2051 ( .A(n308), .B(n309), .S0(next_cr_x[5]), .Y(
        \DP_OP_589J1_125_1438/n25 ) );
  NAND2BXL U2052 ( .AN(n174), .B(next_cr_x[6]), .Y(n309) );
  NAND2XL U2053 ( .A(next_cr_x[6]), .B(n174), .Y(n308) );
  AND2XL U2054 ( .A(next_cr_x[5]), .B(n174), .Y(n230) );
  NAND2XL U2055 ( .A(n1905), .B(n1921), .Y(n1919) );
  NAND2XL U2056 ( .A(n1802), .B(n2712), .Y(n964) );
  INVXL U2057 ( .A(n2710), .Y(n2712) );
  NAND2BXL U2058 ( .AN(n966), .B(n968), .Y(n970) );
  NAND2XL U2059 ( .A(n956), .B(n957), .Y(n955) );
  INVXL U2060 ( .A(n954), .Y(n957) );
  INVXL U2061 ( .A(n959), .Y(n968) );
  INVXL U2062 ( .A(n948), .Y(n952) );
  OAI211XL U2063 ( .A0(write_cntr[1]), .A1(write_cntr[0]), .B0(n946), .C0(n945), .Y(n947) );
  NAND2XL U2064 ( .A(n1803), .B(\intadd_3/A[7] ), .Y(n943) );
  NAND2XL U2065 ( .A(n1021), .B(n1009), .Y(n1020) );
  NAND3XL U2066 ( .A(n1011), .B(n1014), .C(n1012), .Y(n1009) );
  INVXL U2067 ( .A(n1016), .Y(n827) );
  NAND3XL U2068 ( .A(n823), .B(n826), .C(n824), .Y(n822) );
  INVXL U2069 ( .A(n219), .Y(n832) );
  INVXL U2070 ( .A(n843), .Y(n823) );
  INVXL U2071 ( .A(n2717), .Y(\intadd_3/A[7] ) );
  NAND3XL U2072 ( .A(n941), .B(n2754), .C(n940), .Y(n939) );
  NOR2XL U2073 ( .A(n956), .B(n954), .Y(n942) );
  INVXL U2074 ( .A(n953), .Y(n950) );
  NOR2XL U2075 ( .A(n1877), .B(n2761), .Y(n932) );
  NAND2XL U2076 ( .A(n931), .B(n163), .Y(n933) );
  NAND3XL U2077 ( .A(n2750), .B(n2753), .C(n2752), .Y(n2749) );
  AND2XL U2078 ( .A(n2752), .B(n2750), .Y(n2751) );
  NAND2XL U2079 ( .A(n2748), .B(n2747), .Y(n2743) );
  NAND3XL U2080 ( .A(n2748), .B(n2745), .C(n2747), .Y(n2746) );
  NOR2XL U2081 ( .A(n2742), .B(n2741), .Y(n2736) );
  NAND2XL U2082 ( .A(n2742), .B(n2741), .Y(n2739) );
  NAND2XL U2083 ( .A(n2738), .B(n2737), .Y(n2740) );
  NOR2XL U2084 ( .A(n2733), .B(n2731), .Y(n2735) );
  NAND2XL U2085 ( .A(n2722), .B(n2723), .Y(n2721) );
  AND2XL U2086 ( .A(n2720), .B(n226), .Y(n233) );
  OAI31XL U2087 ( .A0(n927), .A1(n161), .A2(n925), .B0(n924), .Y(n934) );
  NOR2BXL U2088 ( .AN(n941), .B(n940), .Y(n928) );
  AND2XL U2089 ( .A(n1880), .B(n2752), .Y(n920) );
  INVXL U2090 ( .A(n935), .Y(n938) );
  NAND2XL U2091 ( .A(n931), .B(n1805), .Y(n935) );
  NAND3XL U2092 ( .A(n161), .B(n922), .C(n923), .Y(n917) );
  OAI31XL U2093 ( .A0(n912), .A1(n911), .A2(n910), .B0(n909), .Y(n926) );
  NOR2XL U2094 ( .A(n907), .B(n906), .Y(n904) );
  NAND2XL U2095 ( .A(n1846), .B(n2737), .Y(n900) );
  NAND2XL U2096 ( .A(n1848), .B(n2730), .Y(n893) );
  NAND2XL U2097 ( .A(n901), .B(n1846), .Y(n902) );
  NOR2XL U2098 ( .A(n896), .B(n897), .Y(n888) );
  INVXL U2099 ( .A(n887), .Y(n890) );
  NAND3XL U2100 ( .A(n881), .B(n2728), .C(n880), .Y(n879) );
  INVXL U2101 ( .A(n878), .Y(n880) );
  NOR2XL U2102 ( .A(n2725), .B(n877), .Y(n875) );
  NAND2BXL U2103 ( .AN(n883), .B(n874), .Y(n876) );
  INVXL U2104 ( .A(n882), .Y(n892) );
  NAND2XL U2105 ( .A(n1848), .B(n894), .Y(n882) );
  NAND2XL U2106 ( .A(n878), .B(n881), .Y(n873) );
  NAND2XL U2107 ( .A(n1806), .B(n2722), .Y(n868) );
  NOR2XL U2108 ( .A(n871), .B(n872), .Y(n862) );
  INVXL U2109 ( .A(n861), .Y(n866) );
  NAND2XL U2110 ( .A(n855), .B(n241), .Y(n854) );
  INVXL U2111 ( .A(n853), .Y(n855) );
  NOR2XL U2112 ( .A(n1018), .B(n2719), .Y(n851) );
  INVXL U2113 ( .A(n856), .Y(n865) );
  NAND2XL U2114 ( .A(n1806), .B(n869), .Y(n856) );
  INVXL U2115 ( .A(n847), .Y(n845) );
  NAND2XL U2116 ( .A(n829), .B(n2718), .Y(n846) );
  NAND2XL U2117 ( .A(n1807), .B(n852), .Y(n850) );
  NOR4XL U2118 ( .A(n809), .B(n808), .C(n812), .D(n945), .Y(n810) );
  NAND2XL U2119 ( .A(write_cntr[1]), .B(write_cntr[0]), .Y(n945) );
  NOR2XL U2120 ( .A(n814), .B(n317), .Y(n813) );
  NAND2XL U2121 ( .A(n829), .B(n847), .Y(n842) );
  AOI211XL U2122 ( .A0(n265), .A1(n815), .B0(n814), .C0(n317), .Y(n840) );
  INVXL U2123 ( .A(n816), .Y(n815) );
  NOR2XL U2124 ( .A(write_cntr[9]), .B(n821), .Y(n820) );
  NAND2XL U2125 ( .A(write_cntr[6]), .B(n837), .Y(n839) );
  NAND4XL U2126 ( .A(write_cntr[5]), .B(write_cntr[3]), .C(write_cntr[2]), .D(
        write_cntr[4]), .Y(n812) );
  INVXL U2127 ( .A(n833), .Y(n834) );
  NAND3XL U2128 ( .A(write_cntr[3]), .B(write_cntr[2]), .C(n930), .Y(n833) );
  NOR2BXL U2129 ( .AN(curr_photo_addr[16]), .B(n313), .Y(\C1/Z_16 ) );
  AOI31XL U2130 ( .A0(n589), .A1(n588), .A2(n587), .B0(n313), .Y(n590) );
  NAND2XL U2131 ( .A(n2832), .B(n586), .Y(n587) );
  INVX3 U2132 ( .A(n740), .Y(\sftr_n[0]_BAR ) );
  NAND2XL U2133 ( .A(n720), .B(\C158/DATA2_16 ), .Y(n588) );
  AOI21XL U2134 ( .A0(n723), .A1(n2830), .B0(n585), .Y(n589) );
  OAI211XL U2135 ( .A0(n710), .A1(n619), .B0(n584), .C0(n583), .Y(n585) );
  NAND2XL U2136 ( .A(n2769), .B(n224), .Y(n365) );
  NOR2BXL U2137 ( .AN(curr_photo_addr[17]), .B(n313), .Y(\C1/Z_17 ) );
  AOI211XL U2138 ( .A0(n2777), .A1(n2776), .B0(n2779), .C0(n2783), .Y(n2778)
         );
  XNOR2XL U2139 ( .A(n366), .B(write_addr[15]), .Y(n367) );
  NAND2BXL U2140 ( .AN(n2769), .B(write_addr[14]), .Y(n366) );
  INVXL U2141 ( .A(n579), .Y(n580) );
  NAND2XL U2142 ( .A(n2806), .B(n2807), .Y(n578) );
  NAND2XL U2143 ( .A(n2802), .B(n2801), .Y(n2808) );
  NAND2XL U2144 ( .A(n2804), .B(n235), .Y(n2801) );
  OAI211XL U2145 ( .A0(n285), .A1(n2804), .B0(n235), .C0(n2799), .Y(n2800) );
  NOR2BXL U2146 ( .AN(curr_photo_addr[18]), .B(n313), .Y(\C1/Z_18 ) );
  AOI211XL U2147 ( .A0(\DP_OP_559J1_134_6328/n1 ), .A1(n720), .B0(n576), .C0(
        n575), .Y(n577) );
  OAI211XL U2148 ( .A0(n603), .A1(n710), .B0(n574), .C0(n573), .Y(n575) );
  NAND2XL U2149 ( .A(n636), .B(write_addr[16]), .Y(n573) );
  INVXL U2150 ( .A(n704), .Y(n636) );
  INVXL U2151 ( .A(n742), .Y(n2794) );
  INVXL U2152 ( .A(n2779), .Y(n2780) );
  NAND2BXL U2153 ( .AN(n2814), .B(n568), .Y(n569) );
  INVXL U2154 ( .A(n567), .Y(n568) );
  AOI211XL U2155 ( .A0(n2872), .A1(n284), .B0(n2873), .C0(n2813), .Y(n2814) );
  INVXL U2156 ( .A(n2771), .Y(n369) );
  INVXL U2157 ( .A(n2772), .Y(n368) );
  AND2XL U2158 ( .A(n2773), .B(n2774), .Y(n2770) );
  OAI211XL U2159 ( .A0(n741), .A1(n2835), .B0(n2838), .C0(n2839), .Y(n1819) );
  NAND2XL U2160 ( .A(write_addr[2]), .B(write_addr[1]), .Y(n1915) );
  INVXL U2161 ( .A(n2840), .Y(n1820) );
  NAND4BXL U2162 ( .AN(n1816), .B(n2775), .C(n2781), .D(n2777), .Y(n1821) );
  NAND2XL U2163 ( .A(write_addr[8]), .B(n2827), .Y(n1815) );
  NAND2XL U2164 ( .A(write_addr[13]), .B(n1811), .Y(n2768) );
  AOI211XL U2165 ( .A0(n2756), .A1(n1810), .B0(n2766), .C0(n1812), .Y(n1816)
         );
  INVXL U2166 ( .A(n2763), .Y(n1810) );
  NOR2XL U2167 ( .A(n223), .B(n1808), .Y(n1809) );
  INVXL U2168 ( .A(n1808), .Y(n2713) );
  INVXL U2169 ( .A(n17), .Y(n1945) );
  OAI31X1 U2170 ( .A0(n27), .A1(n800), .A2(n337), .B0(n799), .Y(next_state[2])
         );
  INVXL U2171 ( .A(n748), .Y(n337) );
  NAND2XL U2172 ( .A(n748), .B(n800), .Y(n802) );
  AOI211XL U2173 ( .A0(n795), .A1(n794), .B0(n793), .C0(n256), .Y(n796) );
  INVXL U2174 ( .A(n757), .Y(n793) );
  OAI211XL U2175 ( .A0(n753), .A1(n792), .B0(n752), .C0(global_cntr[11]), .Y(
        n794) );
  INVXL U2176 ( .A(n746), .Y(n788) );
  INVXL U2177 ( .A(en_so), .Y(n339) );
  NAND2X1 U2178 ( .A(write_cntr[14]), .B(n787), .Y(n306) );
  AOI211XL U2179 ( .A0(n786), .A1(n199), .B0(n805), .C0(n809), .Y(n787) );
  NAND2XL U2180 ( .A(write_cntr[13]), .B(write_cntr[12]), .Y(n809) );
  OAI21X1 U2181 ( .A0(write_cntr[9]), .A1(write_cntr[10]), .B0(write_cntr[11]), 
        .Y(n805) );
  NOR4XL U2182 ( .A(n763), .B(n764), .C(n766), .D(n765), .Y(n784) );
  AOI21X1 U2183 ( .A0(n242), .A1(n319), .B0(n320), .Y(n765) );
  INVXL U2184 ( .A(n332), .Y(n329) );
  INVXL U2185 ( .A(n328), .Y(n330) );
  AOI21X1 U2186 ( .A0(n247), .A1(n332), .B0(n331), .Y(n752) );
  XNOR2X1 U2187 ( .A(n758), .B(global_cntr[17]), .Y(n333) );
  NOR2XL U2188 ( .A(n758), .B(n783), .Y(n780) );
  NAND4XL U2189 ( .A(n1553), .B(global_cntr[16]), .C(global_cntr[14]), .D(n778), .Y(n781) );
  NOR3XL U2190 ( .A(global_cntr[6]), .B(n240), .C(n779), .Y(n778) );
  AND2XL U2191 ( .A(n758), .B(n335), .Y(n336) );
  NOR2X1 U2192 ( .A(n218), .B(n256), .Y(n335) );
  NAND2XL U2193 ( .A(global_cntr[17]), .B(n758), .Y(n334) );
  NOR2X1 U2194 ( .A(n247), .B(n332), .Y(n331) );
  NAND2X1 U2195 ( .A(n767), .B(global_cntr[3]), .Y(n319) );
  AND3XL U2196 ( .A(n740), .B(n2833), .C(write_addr[19]), .Y(n576) );
  AND2XL U2197 ( .A(n2802), .B(n2798), .Y(n2807) );
  INVXL U2198 ( .A(n739), .Y(n2798) );
  NOR2XL U2199 ( .A(n2804), .B(write_addr[8]), .Y(n2795) );
  NOR2XL U2200 ( .A(n2810), .B(n2809), .Y(n2857) );
  NAND2XL U2201 ( .A(write_addr[8]), .B(n2803), .Y(n2809) );
  INVXL U2202 ( .A(n2806), .Y(n2803) );
  NAND4XL U2203 ( .A(write_addr[11]), .B(write_addr[12]), .C(n2796), .D(n282), 
        .Y(n2797) );
  NOR4XL U2204 ( .A(write_addr[16]), .B(n2854), .C(n235), .D(n2824), .Y(n2796)
         );
  AND2XL U2205 ( .A(\C1/Z_7 ), .B(write_addr[9]), .Y(n260) );
  NAND2XL U2206 ( .A(n383), .B(n1550), .Y(n2864) );
  INVXL U2207 ( .A(n1552), .Y(n382) );
  NAND2XL U2208 ( .A(n742), .B(n271), .Y(n565) );
  AOI21X1 U2209 ( .A0(curr_photo_size[0]), .A1(n356), .B0(n1784), .Y(n271) );
  NOR2XL U2210 ( .A(n1547), .B(n1545), .Y(n1546) );
  AND2XL U2211 ( .A(n1544), .B(n284), .Y(n1545) );
  NAND2XL U2212 ( .A(n1543), .B(n1542), .Y(n1547) );
  MXI2XL U2213 ( .A(n1539), .B(n1538), .S0(n1537), .Y(n1540) );
  INVXL U2214 ( .A(n1536), .Y(n1539) );
  AOI21XL U2215 ( .A0(n1544), .A1(n1542), .B0(n284), .Y(n1541) );
  AND2XL U2216 ( .A(n1537), .B(n1538), .Y(n1535) );
  NAND2XL U2217 ( .A(N1825), .B(n1532), .Y(n1544) );
  NOR2XL U2218 ( .A(n1536), .B(n1537), .Y(n1532) );
  NAND2XL U2219 ( .A(n1530), .B(n1533), .Y(n1529) );
  NOR2XL U2220 ( .A(N1826), .B(n1530), .Y(n1526) );
  NAND2XL U2221 ( .A(n1531), .B(n1525), .Y(n1534) );
  INVXL U2222 ( .A(n1520), .Y(n1518) );
  INVXL U2223 ( .A(n1517), .Y(n1522) );
  INVXL U2224 ( .A(n1527), .Y(n1531) );
  NOR2XL U2225 ( .A(N1827), .B(n1517), .Y(n1516) );
  NAND2XL U2226 ( .A(n1515), .B(n1520), .Y(n1524) );
  NAND2XL U2227 ( .A(n1512), .B(n1514), .Y(n1520) );
  NAND2XL U2228 ( .A(n147), .B(n1510), .Y(n1514) );
  NAND2XL U2229 ( .A(n1507), .B(n1506), .Y(n1510) );
  NOR2XL U2230 ( .A(work_cntr[4]), .B(n1500), .Y(n1505) );
  INVXL U2231 ( .A(n1500), .Y(n1509) );
  NAND2XL U2232 ( .A(n1499), .B(n1498), .Y(n1507) );
  NAND2XL U2233 ( .A(n1504), .B(n221), .Y(n1499) );
  NAND2BXL U2234 ( .AN(n1498), .B(n1501), .Y(n1506) );
  NAND2XL U2235 ( .A(n1494), .B(n1493), .Y(n1497) );
  NAND2XL U2236 ( .A(n1492), .B(n1496), .Y(n1491) );
  INVXL U2237 ( .A(n1484), .Y(n1488) );
  NOR2XL U2238 ( .A(work_cntr[6]), .B(n1492), .Y(n1489) );
  INVXL U2239 ( .A(n1485), .Y(n1481) );
  INVXL U2240 ( .A(n1490), .Y(n1493) );
  NOR2XL U2241 ( .A(work_cntr[7]), .B(n1484), .Y(n1479) );
  NAND2XL U2242 ( .A(n1480), .B(n1485), .Y(n1483) );
  NAND2XL U2243 ( .A(n1476), .B(n1478), .Y(n1485) );
  NAND2BXL U2244 ( .AN(n1475), .B(n1474), .Y(n1478) );
  NAND2XL U2245 ( .A(n1471), .B(n1470), .Y(n1474) );
  NAND2XL U2246 ( .A(n1475), .B(n1469), .Y(n1476) );
  NAND2XL U2247 ( .A(n140), .B(n266), .Y(n1469) );
  NAND2XL U2248 ( .A(n1467), .B(n1465), .Y(n1466) );
  NOR2XL U2249 ( .A(work_cntr[9]), .B(n1467), .Y(n1464) );
  NAND2XL U2250 ( .A(n132), .B(n1468), .Y(n1470) );
  NAND2BXL U2251 ( .AN(n1460), .B(n1459), .Y(n1463) );
  NAND2XL U2252 ( .A(n1456), .B(n1455), .Y(n1459) );
  NAND2XL U2253 ( .A(n1460), .B(n1454), .Y(n1461) );
  NAND2XL U2254 ( .A(n1458), .B(n228), .Y(n1454) );
  NAND2XL U2255 ( .A(n1452), .B(n1450), .Y(n1451) );
  NOR2XL U2256 ( .A(work_cntr[11]), .B(n1452), .Y(n1449) );
  NAND2XL U2257 ( .A(n146), .B(n1453), .Y(n1455) );
  NAND2BXL U2258 ( .AN(n1444), .B(n1443), .Y(n1447) );
  NAND2XL U2259 ( .A(n1438), .B(n1444), .Y(n1445) );
  NAND2XL U2260 ( .A(n1436), .B(n1434), .Y(n1435) );
  NAND2XL U2261 ( .A(n1442), .B(n217), .Y(n1438) );
  NOR2XL U2262 ( .A(work_cntr[13]), .B(n1436), .Y(n1432) );
  NAND2XL U2263 ( .A(n1431), .B(n1437), .Y(n1439) );
  INVXL U2264 ( .A(n1433), .Y(n1437) );
  NAND2XL U2265 ( .A(n1427), .B(n1426), .Y(n1430) );
  INVXL U2266 ( .A(n1426), .Y(n1423) );
  NOR2BXL U2267 ( .AN(n1425), .B(work_cntr[14]), .Y(n1419) );
  NAND2XL U2268 ( .A(n227), .B(n1415), .Y(n1417) );
  AND2XL U2269 ( .A(n1418), .B(n227), .Y(n1411) );
  NOR2XL U2270 ( .A(work_cntr[16]), .B(n1410), .Y(n1408) );
  NAND2XL U2271 ( .A(n2812), .B(n2813), .Y(n2868) );
  NAND2XL U2272 ( .A(n2668), .B(n1403), .Y(n1404) );
  INVXL U2273 ( .A(n1644), .Y(n1645) );
  NAND2XL U2274 ( .A(n1952), .B(n1398), .Y(n1399) );
  OAI211XL U2275 ( .A0(n2658), .A1(n1398), .B0(n1397), .C0(n1780), .Y(n1400)
         );
  NAND2XL U2276 ( .A(n1396), .B(n1395), .Y(n1398) );
  NAND2XL U2277 ( .A(n2654), .B(n1394), .Y(n1395) );
  NAND3XL U2278 ( .A(n138), .B(n1393), .C(n2654), .Y(n1391) );
  OAI211XL U2279 ( .A0(n138), .A1(n2654), .B0(n1393), .C0(n1394), .Y(n1392) );
  INVXL U2280 ( .A(n1390), .Y(n1388) );
  NOR2XL U2281 ( .A(n1379), .B(n1383), .Y(n1380) );
  NAND3XL U2282 ( .A(n1373), .B(n1372), .C(n1369), .Y(n1371) );
  INVXL U2283 ( .A(n1368), .Y(n1373) );
  INVXL U2284 ( .A(n1361), .Y(n1363) );
  INVXL U2285 ( .A(n1372), .Y(n1365) );
  NOR2XL U2286 ( .A(n1354), .B(n1353), .Y(n1355) );
  NAND3XL U2287 ( .A(n1359), .B(n1362), .C(n1356), .Y(n1369) );
  NAND3XL U2288 ( .A(n1358), .B(n1357), .C(n1352), .Y(n1356) );
  INVXL U2289 ( .A(n1351), .Y(n1358) );
  NOR2XL U2290 ( .A(n1354), .B(n1723), .Y(n1340) );
  INVXL U2291 ( .A(n1357), .Y(n1349) );
  NOR2XL U2292 ( .A(n1354), .B(n2380), .Y(n1339) );
  NAND3XL U2293 ( .A(n1344), .B(n1338), .C(n1341), .Y(n1352) );
  NAND3XL U2294 ( .A(n1343), .B(n1337), .C(n1342), .Y(n1341) );
  INVXL U2295 ( .A(n1336), .Y(n1342) );
  NAND2XL U2296 ( .A(n1333), .B(n1329), .Y(n1330) );
  NAND2XL U2297 ( .A(n1336), .B(n217), .Y(n1332) );
  INVXL U2298 ( .A(n1338), .Y(n1345) );
  NAND2XL U2299 ( .A(n1402), .B(n1705), .Y(n1327) );
  NAND2BXL U2300 ( .AN(n1331), .B(n1329), .Y(n1337) );
  NAND2BXL U2301 ( .AN(n1333), .B(n1326), .Y(n1331) );
  NAND3XL U2302 ( .A(n1324), .B(n1321), .C(n1323), .Y(n1322) );
  NOR2XL U2303 ( .A(work_cntr[14]), .B(n157), .Y(n1325) );
  INVXL U2304 ( .A(n1323), .Y(n1317) );
  NOR2XL U2305 ( .A(n1354), .B(n1689), .Y(n1311) );
  INVXL U2306 ( .A(n1306), .Y(n1304) );
  NAND2XL U2307 ( .A(n1297), .B(n1296), .Y(n1303) );
  NAND2XL U2308 ( .A(n1300), .B(n1301), .Y(n1295) );
  NOR2XL U2309 ( .A(n1288), .B(n259), .Y(n1291) );
  AOI211XL U2310 ( .A0(work_cntr[19]), .A1(n252), .B0(n1294), .C0(n1285), .Y(
        n1286) );
  NOR2XL U2311 ( .A(n1354), .B(n2379), .Y(n1285) );
  INVXL U2312 ( .A(n1289), .Y(n1294) );
  NAND2XL U2313 ( .A(n1284), .B(work_cntr[17]), .Y(n1289) );
  INVXL U2314 ( .A(n1293), .Y(n1287) );
  NAND2XL U2315 ( .A(n259), .B(n1288), .Y(n1293) );
  INVXL U2316 ( .A(n1299), .Y(n1301) );
  AND2XL U2317 ( .A(n1298), .B(n227), .Y(n1282) );
  INVXL U2318 ( .A(n1310), .Y(n1313) );
  NAND3XL U2319 ( .A(n217), .B(n1402), .C(n2414), .Y(n1310) );
  NOR2XL U2320 ( .A(n1354), .B(n2446), .Y(n1281) );
  INVXL U2321 ( .A(n1730), .Y(n1353) );
  NOR2XL U2322 ( .A(work_cntr[4]), .B(n1354), .Y(n1280) );
  NOR2X1 U2323 ( .A(n378), .B(curr_photo_size[1]), .Y(n379) );
  OAI211XL U2324 ( .A0(n1274), .A1(n1273), .B0(n1272), .C0(n1271), .Y(n1275)
         );
  NAND2BXL U2325 ( .AN(n1276), .B(n1265), .Y(n1273) );
  NAND2XL U2326 ( .A(n1264), .B(n1263), .Y(n1277) );
  INVXL U2327 ( .A(n1265), .Y(n1263) );
  NAND2XL U2328 ( .A(n1251), .B(n1250), .Y(n1276) );
  INVXL U2329 ( .A(n1244), .Y(n1249) );
  INVXL U2330 ( .A(n1242), .Y(n1243) );
  NAND2XL U2331 ( .A(n1239), .B(n1250), .Y(n1242) );
  NOR2BXL U2332 ( .AN(n1247), .B(n1246), .Y(n1239) );
  NOR2XL U2333 ( .A(n1237), .B(n1254), .Y(n1238) );
  NAND2XL U2334 ( .A(n1257), .B(n1256), .Y(n1254) );
  NAND2BXL U2335 ( .AN(n1231), .B(n1230), .Y(n1260) );
  NAND2BXL U2336 ( .AN(n1241), .B(n1240), .Y(n1223) );
  NAND4BXL U2337 ( .AN(n1253), .B(n1219), .C(n232), .D(n1256), .Y(n1225) );
  INVXL U2338 ( .A(n1214), .Y(n1215) );
  INVXL U2339 ( .A(n1250), .Y(n1226) );
  NAND2XL U2340 ( .A(n1210), .B(n1244), .Y(n1211) );
  AND2XL U2341 ( .A(n1235), .B(n1234), .Y(n1245) );
  NOR2XL U2342 ( .A(n1221), .B(n1220), .Y(n1206) );
  NAND2XL U2343 ( .A(n1233), .B(n1235), .Y(n1201) );
  NAND3XL U2344 ( .A(n263), .B(n1218), .C(n1270), .Y(n1209) );
  AND2XL U2345 ( .A(n1176), .B(n1202), .Y(n1177) );
  NAND4XL U2346 ( .A(n1233), .B(n1185), .C(n273), .D(n1187), .Y(n1180) );
  NAND2XL U2347 ( .A(work_cntr[4]), .B(n1164), .Y(n1188) );
  NOR2XL U2348 ( .A(n1168), .B(n1169), .Y(n1162) );
  NAND2XL U2349 ( .A(n1154), .B(n1153), .Y(n1178) );
  INVXL U2350 ( .A(n1175), .Y(n1202) );
  INVXL U2351 ( .A(n1144), .Y(n1146) );
  INVXL U2352 ( .A(n1197), .Y(n1163) );
  NAND2XL U2353 ( .A(n1145), .B(n1144), .Y(n1143) );
  NAND2BXL U2354 ( .AN(n1128), .B(n1127), .Y(n1155) );
  NAND4XL U2355 ( .A(n1152), .B(n1154), .C(n221), .D(n1126), .Y(n1133) );
  NAND2XL U2356 ( .A(n1182), .B(n1183), .Y(n1156) );
  NOR2XL U2357 ( .A(n1119), .B(n1118), .Y(n1120) );
  NAND2XL U2358 ( .A(n1124), .B(n1125), .Y(n1116) );
  NOR2XL U2359 ( .A(n1124), .B(n1125), .Y(n1117) );
  INVXL U2360 ( .A(n1148), .Y(n1134) );
  NAND3XL U2361 ( .A(n172), .B(n1104), .C(n1113), .Y(n1128) );
  OAI2BB2XL U2362 ( .B0(n1103), .B1(n1102), .A0N(n1103), .A1N(n1102), .Y(n1115) );
  NAND2XL U2363 ( .A(n1094), .B(n1096), .Y(n1093) );
  NAND2BXL U2364 ( .AN(n1091), .B(n1095), .Y(n1092) );
  INVXL U2365 ( .A(n1087), .Y(n1090) );
  NOR2BXL U2366 ( .AN(n1094), .B(n1096), .Y(n1091) );
  NAND4XL U2367 ( .A(n1104), .B(n1108), .C(n1097), .D(n268), .Y(n1086) );
  INVXL U2368 ( .A(n1082), .Y(n1083) );
  INVXL U2369 ( .A(n1075), .Y(n1077) );
  INVXL U2370 ( .A(n1106), .Y(n1073) );
  INVXL U2371 ( .A(n1070), .Y(n1069) );
  NAND2XL U2372 ( .A(n1067), .B(n1066), .Y(n1070) );
  NAND2BXL U2373 ( .AN(n1105), .B(n1108), .Y(n1064) );
  NAND2XL U2374 ( .A(n1121), .B(n217), .Y(n1066) );
  NAND2XL U2375 ( .A(n1060), .B(n1085), .Y(n1082) );
  NOR2XL U2376 ( .A(n1051), .B(n1050), .Y(n1054) );
  NAND4XL U2377 ( .A(n1049), .B(n1060), .C(n217), .D(n2423), .Y(n1056) );
  NOR2XL U2378 ( .A(work_cntr[14]), .B(n1046), .Y(n1048) );
  NAND2XL U2379 ( .A(work_cntr[9]), .B(n1045), .Y(n1075) );
  INVXL U2380 ( .A(n1044), .Y(n1076) );
  INVXL U2381 ( .A(n1051), .Y(n1041) );
  NAND2XL U2382 ( .A(n1040), .B(n1044), .Y(n1067) );
  AND2XL U2383 ( .A(n1057), .B(n1053), .Y(n1045) );
  INVXL U2384 ( .A(n1059), .Y(n1053) );
  NAND2XL U2385 ( .A(n1413), .B(n257), .Y(n1412) );
  NAND2XL U2386 ( .A(n1052), .B(n1058), .Y(n1057) );
  NAND4BXL U2387 ( .AN(n1038), .B(n261), .C(n227), .D(n1055), .Y(n1052) );
  INVXL U2388 ( .A(n2515), .Y(n2518) );
  NOR2XL U2389 ( .A(n1283), .B(n2515), .Y(n1037) );
  NAND3XL U2390 ( .A(n1040), .B(n1068), .C(n1049), .Y(n1038) );
  INVXL U2391 ( .A(n1061), .Y(n1071) );
  INVXL U2392 ( .A(n1035), .Y(n1046) );
  INVXL U2393 ( .A(n1043), .Y(n1034) );
  NAND2XL U2394 ( .A(work_cntr[10]), .B(n1036), .Y(n1042) );
  NAND3XL U2395 ( .A(write_cntr[8]), .B(write_cntr[10]), .C(n1588), .Y(n1562)
         );
  OAI31XL U2396 ( .A0(n2868), .A1(n2867), .A2(n2866), .B0(n2865), .Y(n2869) );
  AOI211XL U2397 ( .A0(n2675), .A1(n2674), .B0(curr_photo_size[0]), .C0(n2673), 
        .Y(n2676) );
  OAI211XL U2398 ( .A0(n1787), .A1(n1786), .B0(curr_photo_size[0]), .C0(n775), 
        .Y(n1795) );
  NAND2BXL U2399 ( .AN(n1549), .B(curr_photo_size[1]), .Y(n356) );
  OAI22XL U2400 ( .A0(n2793), .A1(n381), .B0(n2792), .B1(n304), .Y(
        next_photo[1]) );
  OR2X1 U2401 ( .A(n1636), .B(n385), .Y(n424) );
  NAND3XL U2402 ( .A(write_cntr[9]), .B(write_cntr[11]), .C(write_cntr[10]), 
        .Y(n1558) );
  NOR2XL U2403 ( .A(N196), .B(n232), .Y(n1641) );
  NAND2X1 U2404 ( .A(n318), .B(n2875), .Y(so_mux_sel[1]) );
  NAND2XL U2405 ( .A(N196), .B(n232), .Y(n2861) );
  OAI22XL U2406 ( .A0(n2876), .A1(n237), .B0(n2877), .B1(n2811), .Y(n472) );
  MXI2XL U2407 ( .A(n2699), .B(n2690), .S0(N1138), .Y(n454) );
  AOI21XL U2408 ( .A0(n2695), .A1(N1138), .B0(N1139), .Y(n380) );
  OAI22XL U2409 ( .A0(n2692), .A1(n2691), .B0(n2690), .B1(n302), .Y(n450) );
  OAI2BB2XL U2410 ( .B0(n2703), .B1(n2702), .A0N(cr_read_cntr[8]), .A1N(n2701), 
        .Y(n446) );
  OAI22XL U2411 ( .A0(n224), .A1(n2785), .B0(im_wen_n), .B1(n619), .Y(n439) );
  OAI22XL U2412 ( .A0(n135), .A1(n283), .B0(im_wen_n), .B1(n158), .Y(n436) );
  OAI22XL U2413 ( .A0(n134), .A1(n1804), .B0(n2785), .B1(n269), .Y(n497) );
  OAI21XL U2414 ( .A0(n603), .A1(n134), .B0(n372), .Y(n437) );
  OAI21XL U2415 ( .A0(n134), .A1(n716), .B0(n377), .Y(n482) );
  OAI21XL U2416 ( .A0(n134), .A1(n675), .B0(n361), .Y(n477) );
  OAI21XL U2417 ( .A0(n238), .A1(n135), .B0(n357), .Y(n480) );
  OAI21XL U2418 ( .A0(n2846), .A1(n134), .B0(n374), .Y(n445) );
  OAI22XL U2419 ( .A0(n281), .A1(n135), .B0(im_wen_n), .B1(n373), .Y(n435) );
  OAI2BB2XL U2420 ( .B0(n134), .B1(n1803), .A0N(n134), .A1N(write_cntr[2]), 
        .Y(n499) );
  OAI22XL U2421 ( .A0(n282), .A1(n135), .B0(im_wen_n), .B1(n375), .Y(n434) );
  OAI22XL U2422 ( .A0(n299), .A1(n135), .B0(im_wen_n), .B1(n607), .Y(n438) );
  OAI21XL U2423 ( .A0(n134), .A1(n701), .B0(n359), .Y(n479) );
  OAI21XL U2424 ( .A0(n134), .A1(n2852), .B0(n363), .Y(n475) );
  OAI22XL U2425 ( .A0(n134), .A1(n219), .B0(n135), .B1(n234), .Y(n485) );
  OAI22XL U2426 ( .A0(n134), .A1(n1807), .B0(n135), .B1(n199), .Y(n489) );
  OAI22XL U2427 ( .A0(n134), .A1(n1897), .B0(n135), .B1(n220), .Y(n495) );
  OAI22XL U2428 ( .A0(n134), .A1(n1848), .B0(n135), .B1(n272), .Y(n491) );
  OAI22XL U2429 ( .A0(n134), .A1(n1846), .B0(n135), .B1(n287), .Y(n492) );
  OAI22XL U2430 ( .A0(n134), .A1(n829), .B0(n135), .B1(n278), .Y(n488) );
  OAI22XL U2431 ( .A0(n134), .A1(n847), .B0(n135), .B1(n265), .Y(n487) );
  OAI22XL U2432 ( .A0(n134), .A1(n1806), .B0(n135), .B1(n267), .Y(n490) );
  OAI22XL U2433 ( .A0(n134), .A1(n1855), .B0(n135), .B1(n274), .Y(n493) );
  OAI22XL U2434 ( .A0(n134), .A1(n841), .B0(n135), .B1(n279), .Y(n486) );
  OAI22XL U2435 ( .A0(n134), .A1(n1880), .B0(n135), .B1(n275), .Y(n498) );
  OAI22XL U2436 ( .A0(n134), .A1(n1805), .B0(n135), .B1(n276), .Y(n494) );
  OAI22XL U2437 ( .A0(n134), .A1(n1802), .B0(n135), .B1(n262), .Y(n500) );
  CLKBUFX3 U2438 ( .A(n728), .Y(n311) );
  OA22X1 U2439 ( .A0(n961), .A1(n811), .B0(n234), .B1(n960), .Y(n219) );
  OR2X1 U2440 ( .A(n2684), .B(n1917), .Y(n2682) );
  CLKBUFX3 U2441 ( .A(n745), .Y(n310) );
  NOR3XL U2442 ( .A(write_cntr[14]), .B(write_cntr[13]), .C(write_cntr[12]), 
        .Y(n806) );
  NAND4XL U2443 ( .A(write_cntr[11]), .B(write_cntr[8]), .C(write_cntr[7]), 
        .D(write_cntr[6]), .Y(n808) );
  CLKBUFX3 U2444 ( .A(si_sel), .Y(n312) );
  AND2X2 U2445 ( .A(n316), .B(n2709), .Y(n744) );
  NOR2X1 U2446 ( .A(n1947), .B(n1945), .Y(n2709) );
  NAND2X1 U2447 ( .A(n804), .B(n803), .Y(n17) );
  NAND3X1 U2448 ( .A(n798), .B(n797), .C(n802), .Y(n804) );
  NOR3X1 U2449 ( .A(n750), .B(n749), .C(n796), .Y(n800) );
  AOI211X1 U2450 ( .A0(n747), .A1(n2681), .B0(n791), .C0(n790), .Y(n798) );
  OAI22XL U2451 ( .A0(n797), .A1(n2111), .B0(n1783), .B1(n801), .Y(n790) );
  AOI221XL U2452 ( .A0(n769), .A1(n1946), .B0(n254), .B1(n1946), .C0(n788), 
        .Y(n791) );
  OAI31XL U2453 ( .A0(write_cntr[7]), .A1(write_cntr[5]), .A2(write_cntr[6]), 
        .B0(write_cntr[8]), .Y(n786) );
  OA21XL U2454 ( .A0(global_cntr[7]), .A1(n326), .B0(n327), .Y(n755) );
  NOR2X1 U2455 ( .A(n783), .B(n333), .Y(n751) );
  OA22X1 U2456 ( .A0(n336), .A1(global_cntr[19]), .B0(n780), .B1(n779), .Y(
        n749) );
  NAND2XL U2457 ( .A(global_cntr[19]), .B(n335), .Y(n779) );
  NOR2X1 U2458 ( .A(n249), .B(n321), .Y(n322) );
  NAND2X1 U2459 ( .A(global_cntr[11]), .B(n331), .Y(n321) );
  NOR2X1 U2460 ( .A(n243), .B(n327), .Y(n328) );
  AND2X2 U2461 ( .A(n769), .B(global_cntr[2]), .Y(n767) );
  INVX3 U2462 ( .A(n314), .Y(n313) );
  INVX3 U2463 ( .A(n725), .Y(n314) );
  CLKINVX1 U2464 ( .A(n1354), .Y(n1402) );
  MXI2X1 U2465 ( .A(n632), .B(n297), .S0(n134), .Y(n441) );
  MXI2X1 U2466 ( .A(n650), .B(n294), .S0(n134), .Y(n444) );
  AOI21X1 U2467 ( .A0(n249), .A1(n321), .B0(n322), .Y(n762) );
  NAND2X1 U2468 ( .A(global_cntr[15]), .B(n324), .Y(n325) );
  NOR2X1 U2469 ( .A(n248), .B(n323), .Y(n324) );
  AOI2BB1X1 U2470 ( .A0N(global_cntr[1]), .A1N(global_cntr[0]), .B0(n769), .Y(
        \next_glb_cntr[1] ) );
  OAI21XL U2471 ( .A0(n469), .A1(n471), .B0(n508), .Y(n470) );
  OAI22XL U2472 ( .A0(n992), .A1(n420), .B0(n993), .B1(n421), .Y(n422) );
  AOI2BB2X1 U2473 ( .B0(n505), .B1(m_1[3]), .A0N(n408), .A1N(n554), .Y(n496)
         );
  OAI22XL U2474 ( .A0(n515), .A1(n528), .B0(n514), .B1(n525), .Y(n516) );
  OAI22XL U2475 ( .A0(n520), .A1(n508), .B0(n507), .B1(n506), .Y(n517) );
  AO21X1 U2476 ( .A0(n503), .A1(n502), .B0(n501), .Y(n504) );
  OR2X1 U2477 ( .A(n533), .B(curr_time[9]), .Y(n502) );
  OAI22XL U2478 ( .A0(n528), .A1(n527), .B0(n526), .B1(n525), .Y(n529) );
  OAI21XL U2479 ( .A0(cr_read_cntr[3]), .A1(n560), .B0(n559), .Y(N89) );
  AO22X1 U2480 ( .A0(n551), .A1(\s_0[0] ), .B0(n550), .B1(n541), .Y(n542) );
  AOI2BB2X1 U2481 ( .B0(n455), .B1(n976), .A0N(n975), .A1N(n457), .Y(n463) );
  AOI2BB2X1 U2482 ( .B0(n456), .B1(n431), .A0N(n973), .A1N(n427), .Y(n428) );
  OR2X1 U2483 ( .A(n1797), .B(n1800), .Y(n547) );
  AOI2BB2X1 U2484 ( .B0(n540), .B1(\m_0[0] ), .A0N(n539), .A1N(n555), .Y(n544)
         );
  OR2X1 U2485 ( .A(n549), .B(n743), .Y(n555) );
  OAI2BB1X1 U2486 ( .A0N(n395), .A1N(n394), .B0(n392), .Y(n405) );
  OAI2BB1X1 U2487 ( .A0N(n981), .A1N(n391), .B0(n390), .Y(n396) );
  OR2X1 U2488 ( .A(n387), .B(n386), .Y(n401) );
  AOI2BB1X1 U2489 ( .A0N(n1637), .A1N(n1638), .B0(n1623), .Y(n385) );
  AOI2BB1X1 U2490 ( .A0N(n564), .A1N(n563), .B0(n562), .Y(N88) );
  NAND3BX1 U2491 ( .AN(n1028), .B(n239), .C(n302), .Y(n557) );
  OAI2BB1X1 U2492 ( .A0N(cr_read_cntr[3]), .A1N(n2694), .B0(n2688), .Y(n451)
         );
  NOR2XL U2493 ( .A(n2686), .B(n303), .Y(n2687) );
  OAI211XL U2494 ( .A0(n2506), .A1(n232), .B0(n2507), .C0(n263), .Y(n2505) );
  AOI2BB1X1 U2495 ( .A0N(global_cntr[2]), .A1N(n769), .B0(n767), .Y(n768) );
  NAND2XL U2496 ( .A(n232), .B(n263), .Y(n2497) );
  AO22X1 U2497 ( .A0(n724), .A1(global_cntr[19]), .B0(n314), .B1(n572), .Y(
        \C2/Z_19 ) );
  OR2X1 U2498 ( .A(n704), .B(n283), .Y(n570) );
  AOI2BB2X1 U2499 ( .B0(n582), .B1(n697), .A0N(n718), .A1N(n282), .Y(n571) );
  OAI22XL U2500 ( .A0(n313), .A1(n714), .B0(n1783), .B1(n290), .Y(\C2/Z_1 ) );
  OAI22XL U2501 ( .A0(n704), .A1(n236), .B0(n718), .B1(n288), .Y(n705) );
  AO22X1 U2502 ( .A0(curr_photo_addr[1]), .A1(n314), .B0(n724), .B1(
        curr_photo[0]), .Y(n730) );
  AO22X1 U2503 ( .A0(curr_photo_addr[2]), .A1(n314), .B0(n724), .B1(
        curr_photo[1]), .Y(n731) );
  AO22X1 U2504 ( .A0(n314), .A1(n702), .B0(n724), .B1(global_cntr[2]), .Y(
        \C2/Z_2 ) );
  OAI21XL U2505 ( .A0(n717), .A1(n2835), .B0(n693), .Y(n694) );
  OAI22XL U2506 ( .A0(n704), .A1(n288), .B0(n718), .B1(n238), .Y(n692) );
  OAI2BB1X1 U2507 ( .A0N(curr_photo_addr[3]), .A1N(n314), .B0(n318), .Y(n732)
         );
  OAI22XL U2508 ( .A0(n313), .A1(n691), .B0(n1783), .B1(n291), .Y(\C2/Z_3 ) );
  OAI22XL U2509 ( .A0(n704), .A1(n238), .B0(n718), .B1(n289), .Y(n684) );
  OAI2BB1X1 U2510 ( .A0N(curr_photo_addr[4]), .A1N(n314), .B0(n318), .Y(n733)
         );
  OAI22XL U2511 ( .A0(n313), .A1(n682), .B0(n1783), .B1(n242), .Y(\C2/Z_4 ) );
  OAI22XL U2512 ( .A0(n704), .A1(n289), .B0(n718), .B1(n741), .Y(n676) );
  AO22X1 U2513 ( .A0(n314), .A1(n674), .B0(n724), .B1(global_cntr[5]), .Y(
        \C2/Z_5 ) );
  OAI21XL U2514 ( .A0(n2845), .A1(n700), .B0(n673), .Y(n674) );
  OAI22XL U2515 ( .A0(n704), .A1(n741), .B0(n718), .B1(n293), .Y(n668) );
  AO21X1 U2516 ( .A0(n310), .A1(\intadd_3/SUM[1] ), .B0(n360), .Y(n690) );
  OAI22XL U2517 ( .A0(n683), .A1(n776), .B0(n2771), .B1(n741), .Y(n360) );
  OAI22XL U2518 ( .A0(n313), .A1(n667), .B0(n1783), .B1(n244), .Y(\C2/Z_6 ) );
  OAI22XL U2519 ( .A0(n704), .A1(n293), .B0(n718), .B1(n222), .Y(n660) );
  OAI2BB1X1 U2520 ( .A0N(curr_photo_addr[7]), .A1N(n314), .B0(n318), .Y(n736)
         );
  OAI22XL U2521 ( .A0(n725), .A1(n659), .B0(n1783), .B1(n298), .Y(\C2/Z_7 ) );
  OAI21XL U2522 ( .A0(n2845), .A1(n710), .B0(n656), .Y(n657) );
  OAI31XL U2523 ( .A0(n2844), .A1(\sftr_n[0]_BAR ), .A2(n294), .B0(n653), .Y(
        n654) );
  AOI2BB2X1 U2524 ( .B0(n652), .B1(write_addr[7]), .A0N(n704), .A1N(n222), .Y(
        n653) );
  OAI22XL U2525 ( .A0(n725), .A1(n649), .B0(n1783), .B1(n243), .Y(\C2/Z_8 ) );
  OAI22XL U2526 ( .A0(n704), .A1(n295), .B0(n718), .B1(n235), .Y(n642) );
  OAI22XL U2527 ( .A0(n725), .A1(n641), .B0(n1783), .B1(n247), .Y(\C2/Z_10 )
         );
  OAI31XL U2528 ( .A0(\sftr_n[0]_BAR ), .A1(n2819), .A2(n297), .B0(n633), .Y(
        n634) );
  OAI2BB1X1 U2529 ( .A0N(curr_photo_addr[11]), .A1N(n314), .B0(n318), .Y(
        \C1/Z_11 ) );
  OAI22XL U2530 ( .A0(n725), .A1(n631), .B0(n1783), .B1(n300), .Y(\C2/Z_11 )
         );
  OAI21XL U2531 ( .A0(n650), .A1(n710), .B0(n628), .Y(n629) );
  OAI22XL U2532 ( .A0(n704), .A1(n294), .B0(n718), .B1(n223), .Y(n626) );
  OAI31XL U2533 ( .A0(n2715), .A1(write_addr[9]), .A2(n2711), .B0(n2714), .Y(
        n364) );
  AO22X1 U2534 ( .A0(n314), .A1(n623), .B0(n724), .B1(global_cntr[12]), .Y(
        \C2/Z_12 ) );
  OAI21XL U2535 ( .A0(n632), .A1(n715), .B0(n622), .Y(n623) );
  OAI21XL U2536 ( .A0(n2823), .A1(n296), .B0(n224), .Y(n616) );
  AOI2BB2X1 U2537 ( .B0(n652), .B1(write_addr[12]), .A0N(n704), .A1N(n292), 
        .Y(n618) );
  OAI2BB1X1 U2538 ( .A0N(curr_photo_addr[13]), .A1N(n314), .B0(n318), .Y(
        \C1/Z_13 ) );
  AO22X1 U2539 ( .A0(n314), .A1(n615), .B0(n724), .B1(global_cntr[13]), .Y(
        \C2/Z_13 ) );
  AO21X1 U2540 ( .A0(n2826), .A1(n2822), .B0(write_addr[15]), .Y(n608) );
  OAI2BB1X1 U2541 ( .A0N(curr_photo_addr[14]), .A1N(n314), .B0(n318), .Y(
        \C1/Z_14 ) );
  OAI22XL U2542 ( .A0(n725), .A1(n606), .B0(n1783), .B1(n248), .Y(\C2/Z_14 )
         );
  AOI2BB1X1 U2543 ( .A0N(n704), .A1N(n297), .B0(n599), .Y(n602) );
  OAI22XL U2544 ( .A0(n715), .A1(n619), .B0(n224), .B1(n718), .Y(n599) );
  OAI2BB1X1 U2545 ( .A0N(curr_photo_addr[15]), .A1N(n314), .B0(n318), .Y(
        \C1/Z_15 ) );
  AO22X1 U2546 ( .A0(n314), .A1(n598), .B0(n724), .B1(global_cntr[15]), .Y(
        \C2/Z_15 ) );
  AO21X1 U2547 ( .A0(n2827), .A1(n2826), .B0(write_addr[17]), .Y(n591) );
  AOI31XL U2548 ( .A0(write_cntr[9]), .A1(write_cntr[10]), .A2(n810), .B0(
        write_cntr[14]), .Y(n811) );
  AO21X1 U2549 ( .A0(global_cntr[16]), .A1(n724), .B0(n590), .Y(\C2/Z_16 ) );
  OAI22XL U2550 ( .A0(n717), .A1(n2829), .B0(\sftr_n[0]_BAR ), .B1(n281), .Y(
        n586) );
  OR2X1 U2551 ( .A(n704), .B(n224), .Y(n583) );
  AOI2BB2X1 U2552 ( .B0(n652), .B1(write_addr[16]), .A0N(n603), .A1N(n715), 
        .Y(n584) );
  OAI2BB1X1 U2553 ( .A0N(n285), .A1N(n2808), .B0(n580), .Y(n581) );
  OAI2BB1X1 U2554 ( .A0N(n2810), .A1N(n2805), .B0(n578), .Y(n579) );
  OAI22XL U2555 ( .A0(n313), .A1(n577), .B0(n1783), .B1(n218), .Y(\C2/Z_18 )
         );
  AOI2BB2X1 U2556 ( .B0(n2830), .B1(n697), .A0N(n718), .A1N(n281), .Y(n574) );
  NAND3BX1 U2557 ( .AN(n2815), .B(n285), .C(n237), .Y(n567) );
  OA21XL U2558 ( .A0(global_cntr[13]), .A1(n322), .B0(n323), .Y(n761) );
  OA21XL U2559 ( .A0(global_cntr[15]), .A1(n324), .B0(n325), .Y(n759) );
  OA21XL U2560 ( .A0(global_cntr[3]), .A1(n767), .B0(n319), .Y(n766) );
  OA21XL U2561 ( .A0(global_cntr[5]), .A1(n320), .B0(n782), .Y(n764) );
  OA21XL U2562 ( .A0(global_cntr[11]), .A1(n331), .B0(n321), .Y(n763) );
  AO21X1 U2563 ( .A0(read_cntr[0]), .A1(n739), .B0(n738), .Y(\C1/Z_7 ) );
  OAI2BB1X1 U2564 ( .A0N(n1557), .A1N(n1556), .B0(n384), .Y(n2802) );
  NAND3BX1 U2565 ( .AN(n1551), .B(n284), .C(n382), .Y(n383) );
  OR2X1 U2566 ( .A(n849), .B(n219), .Y(n226) );
  OR2X1 U2567 ( .A(n1030), .B(n1029), .Y(n239) );
  OR2X1 U2568 ( .A(curr_photo_size[0]), .B(n2794), .Y(n286) );
  OR4X1 U2569 ( .A(global_cntr[10]), .B(global_cntr[11]), .C(global_cntr[12]), 
        .D(global_cntr[13]), .Y(n777) );
  CLKINVX1 U2570 ( .A(n789), .Y(n797) );
  OA21XL U2571 ( .A0(n755), .A1(n756), .B0(n754), .Y(n792) );
  OAI22XL U2572 ( .A0(n267), .A1(n817), .B0(n199), .B1(n317), .Y(n818) );
  AOI2BB2X1 U2573 ( .B0(n826), .B1(n825), .A0N(n826), .A1N(n825), .Y(n1011) );
  OAI21XL U2574 ( .A0(n226), .A1(n849), .B0(n219), .Y(n848) );
  OAI21XL U2575 ( .A0(n860), .A1(n857), .B0(n859), .Y(n858) );
  OAI21XL U2576 ( .A0(n865), .A1(n2724), .B0(n864), .Y(n863) );
  OAI21XL U2577 ( .A0(n866), .A1(n1015), .B0(n869), .Y(n867) );
  OAI21XL U2578 ( .A0(n2724), .A1(n871), .B0(n872), .Y(n870) );
  OAI21XL U2579 ( .A0(n886), .A1(n883), .B0(n885), .Y(n884) );
  OAI21XL U2580 ( .A0(n892), .A1(n2733), .B0(n891), .Y(n889) );
  AOI2BB2X1 U2581 ( .B0(n1848), .B1(n2730), .A0N(n1848), .A1N(n2730), .Y(n901)
         );
  OAI21XL U2582 ( .A0(n2733), .A1(n896), .B0(n897), .Y(n895) );
  OAI21XL U2583 ( .A0(n898), .A1(n1857), .B0(n901), .Y(n899) );
  OR2X1 U2584 ( .A(n916), .B(n915), .Y(n908) );
  OAI21XL U2585 ( .A0(n912), .A1(n2744), .B0(n911), .Y(n909) );
  AOI2BB2X1 U2586 ( .B0(n1873), .B1(n2744), .A0N(n1873), .A1N(n2744), .Y(n921)
         );
  OAI21XL U2587 ( .A0(n2744), .A1(n915), .B0(n916), .Y(n914) );
  AOI2BB2X1 U2588 ( .B0(n1880), .B1(n2752), .A0N(n1880), .A1N(n2752), .Y(n931)
         );
  NAND3BX1 U2589 ( .AN(n918), .B(n921), .C(n1880), .Y(n919) );
  AOI2BB2X1 U2590 ( .B0(n923), .B1(n925), .A0N(n923), .A1N(n925), .Y(n940) );
  OAI2BB1X1 U2591 ( .A0N(n923), .A1N(n922), .B0(n161), .Y(n924) );
  OAI2BB1X1 U2592 ( .A0N(n935), .A1N(n163), .B0(n937), .Y(n936) );
  AOI2BB2X1 U2593 ( .B0(n2717), .B1(n1803), .A0N(n2717), .A1N(n1803), .Y(n965)
         );
  OAI2BB1X1 U2594 ( .A0N(n950), .A1N(n949), .B0(n952), .Y(n951) );
  OAI2BB1X1 U2595 ( .A0N(n968), .A1N(n969), .B0(n963), .Y(n958) );
  AOI2BB2X1 U2596 ( .B0(n1802), .B1(n2710), .A0N(n1802), .A1N(n2710), .Y(n1900) );
  OA22X1 U2597 ( .A0(n970), .A1(n2710), .B0(n969), .B1(n968), .Y(n1921) );
  OR2X1 U2598 ( .A(n976), .B(curr_time[19]), .Y(n975) );
  AOI2BB2X1 U2599 ( .B0(n995), .B1(n231), .A0N(n995), .A1N(n231), .Y(n2519) );
  AOI2BB2X1 U2600 ( .B0(n1014), .B1(n1013), .A0N(n1014), .A1N(n1013), .Y(n1828) );
  AOI2BB2X1 U2601 ( .B0(n1031), .B1(n1030), .A0N(n1031), .A1N(n1030), .Y(n1033) );
  NAND3BX1 U2602 ( .AN(n1642), .B(n216), .C(n227), .Y(n1039) );
  OA22X1 U2603 ( .A0(n1037), .A1(n231), .B0(n1283), .B1(n1407), .Y(n1055) );
  AOI2BB1X1 U2604 ( .A0N(n1283), .A1N(n1407), .B0(n252), .Y(n1058) );
  AOI2BB2X1 U2605 ( .B0(n1050), .B1(n1041), .A0N(n1050), .A1N(n1041), .Y(n1065) );
  OAI21XL U2606 ( .A0(n1081), .A1(work_cntr[11]), .B0(work_cntr[12]), .Y(n1080) );
  OR2X1 U2607 ( .A(n1142), .B(n1174), .Y(n1138) );
  AOI2BB2X1 U2608 ( .B0(n1123), .B1(n1122), .A0N(n1123), .A1N(n1122), .Y(n1183) );
  AOI2BB2X1 U2609 ( .B0(n1132), .B1(n1131), .A0N(n1132), .A1N(n1131), .Y(n1147) );
  OAI21XL U2610 ( .A0(n1151), .A1(n1153), .B0(n1154), .Y(n1150) );
  AND4X1 U2611 ( .A(n270), .B(n1202), .C(n1152), .D(n1160), .Y(n1159) );
  OA21XL U2612 ( .A0(n1156), .A1(n1178), .B0(n1155), .Y(n1157) );
  AOI2BB2X1 U2613 ( .B0(n1158), .B1(n1157), .A0N(n1158), .A1N(n1157), .Y(n1167) );
  AO21X1 U2614 ( .A0(n1167), .A1(n1166), .B0(n1165), .Y(n1205) );
  NAND4BBXL U2615 ( .AN(n1180), .BN(n1221), .C(n1207), .D(n1203), .Y(n1204) );
  AOI2BB2X1 U2616 ( .B0(n1184), .B1(n1183), .A0N(n1184), .A1N(n1183), .Y(n1195) );
  NAND4BBXL U2617 ( .AN(n1222), .BN(n1209), .C(n1219), .D(n1202), .Y(n1208) );
  AOI2BB2X1 U2618 ( .B0(n1218), .B1(n1217), .A0N(n1218), .A1N(n1217), .Y(n1256) );
  AOI2BB2X1 U2619 ( .B0(n1221), .B1(n1220), .A0N(n1221), .A1N(n1220), .Y(n1224) );
  AOI2BB2X1 U2620 ( .B0(n1224), .B1(n1223), .A0N(n1224), .A1N(n1223), .Y(n1231) );
  OAI21XL U2621 ( .A0(n1247), .A1(n1245), .B0(n1246), .Y(n1248) );
  OAI22XL U2622 ( .A0(n1249), .A1(n1248), .B0(n1247), .B1(n1246), .Y(n1251) );
  NOR3BXL U2623 ( .AN(n1254), .B(n1253), .C(n1252), .Y(n1255) );
  OA21XL U2624 ( .A0(n1257), .A1(n1256), .B0(n1255), .Y(n1272) );
  NAND3BX1 U2625 ( .AN(n1276), .B(n1272), .C(n1265), .Y(n1259) );
  AOI2BB2X1 U2626 ( .B0(n1270), .B1(n1269), .A0N(n1270), .A1N(n1269), .Y(n1271) );
  AOI2BB1X1 U2627 ( .A0N(n1354), .A1N(n2379), .B0(n252), .Y(n1288) );
  OAI21XL U2628 ( .A0(n2379), .A1(n1354), .B0(n1289), .Y(n1290) );
  NAND3BX1 U2629 ( .AN(n1292), .B(n1291), .C(n1290), .Y(n1296) );
  AOI222XL U2630 ( .A0(n1300), .A1(n1308), .B0(n1300), .B1(work_cntr[16]), 
        .C0(n1308), .C1(n1299), .Y(n1302) );
  AOI2BB2X1 U2631 ( .B0(n1303), .B1(n1302), .A0N(n1303), .A1N(n1301), .Y(n1307) );
  OAI21XL U2632 ( .A0(work_cntr[15]), .A1(n1316), .B0(n1307), .Y(n1305) );
  AOI2BB2X1 U2633 ( .B0(n1308), .B1(n1307), .A0N(n1308), .A1N(n1307), .Y(n1320) );
  OAI21XL U2634 ( .A0(n157), .A1(n1314), .B0(n1316), .Y(n1309) );
  OR2X1 U2635 ( .A(n1314), .B(n157), .Y(n1315) );
  OAI2BB1X1 U2636 ( .A0N(n1316), .A1N(n157), .B0(n1315), .Y(n1323) );
  OAI31XL U2637 ( .A0(n1324), .A1(work_cntr[14]), .A2(n157), .B0(n1317), .Y(
        n1318) );
  AOI2BB1X1 U2638 ( .A0N(work_cntr[13]), .A1N(n1329), .B0(n1318), .Y(n1319) );
  AOI2BB2X1 U2639 ( .B0(n1321), .B1(n1319), .A0N(n1321), .A1N(n1324), .Y(n1326) );
  OA21XL U2640 ( .A0(n1326), .A1(n1329), .B0(n1337), .Y(n1335) );
  AO21X1 U2641 ( .A0(n251), .A1(n1345), .B0(n1343), .Y(n1334) );
  OA21XL U2642 ( .A0(n1344), .A1(n1338), .B0(n1352), .Y(n1350) );
  AO21X1 U2643 ( .A0(n228), .A1(n1349), .B0(n1344), .Y(n1346) );
  OAI21XL U2644 ( .A0(work_cntr[9]), .A1(n1362), .B0(n1351), .Y(n1348) );
  AO21X1 U2645 ( .A0(n266), .A1(n1365), .B0(n1359), .Y(n1360) );
  OAI21XL U2646 ( .A0(work_cntr[7]), .A1(n1367), .B0(n1368), .Y(n1364) );
  AOI2BB2X1 U2647 ( .B0(n1366), .B1(n1365), .A0N(n1366), .A1N(n1364), .Y(n1370) );
  OA21XL U2648 ( .A0(n1373), .A1(n1372), .B0(n1371), .Y(n1377) );
  OAI21XL U2649 ( .A0(work_cntr[6]), .A1(n1386), .B0(n1374), .Y(n1376) );
  OAI21XL U2650 ( .A0(work_cntr[5]), .A1(n1387), .B0(n1385), .Y(n1378) );
  NOR3BXL U2651 ( .AN(n1386), .B(n1383), .C(n1385), .Y(n1381) );
  OAI21XL U2652 ( .A0(n1383), .A1(n1385), .B0(n1386), .Y(n1384) );
  AO21X1 U2653 ( .A0(n2654), .A1(n1393), .B0(n1394), .Y(n1396) );
  AOI2BB2X1 U2654 ( .B0(n1405), .B1(n1400), .A0N(n1405), .A1N(n1399), .Y(n1403) );
  AOI2BB2X1 U2655 ( .B0(n2668), .B1(n1403), .A0N(n2668), .A1N(n1403), .Y(n2872) );
  AOI2BB2X1 U2656 ( .B0(n1405), .B1(n1404), .A0N(n1405), .A1N(n1404), .Y(n1406) );
  AOI2BB2X1 U2657 ( .B0(n1406), .B1(n2658), .A0N(n1406), .A1N(n2658), .Y(n2813) );
  OAI22XL U2658 ( .A0(n2862), .A1(n2868), .B0(n2496), .B1(n2812), .Y(n1549) );
  OA21XL U2659 ( .A0(work_cntr[19]), .A1(n231), .B0(n1407), .Y(n1409) );
  OR2X1 U2660 ( .A(n1409), .B(n1408), .Y(n1422) );
  AO21X1 U2661 ( .A0(n1412), .A1(n1422), .B0(n1411), .Y(n1420) );
  AOI2BB1X1 U2662 ( .A0N(n252), .A1N(n1414), .B0(n1413), .Y(n1421) );
  AOI2BB2X1 U2663 ( .B0(n227), .B1(n1415), .A0N(n227), .A1N(n1415), .Y(n1425)
         );
  OAI21XL U2664 ( .A0(work_cntr[15]), .A1(n1421), .B0(n1418), .Y(n1416) );
  OAI2BB1X1 U2665 ( .A0N(n1422), .A1N(n1421), .B0(n1420), .Y(n1426) );
  OAI21XL U2666 ( .A0(n1426), .A1(work_cntr[14]), .B0(n1425), .Y(n1424) );
  OA21XL U2667 ( .A0(n2423), .A1(n1439), .B0(n1434), .Y(n1442) );
  OAI2BB1X1 U2668 ( .A0N(n1445), .A1N(n1443), .B0(n217), .Y(n1446) );
  OAI21XL U2669 ( .A0(n1443), .A1(work_cntr[12]), .B0(n1442), .Y(n1441) );
  OR2X1 U2670 ( .A(n1449), .B(n146), .Y(n1456) );
  OAI2BB1X1 U2671 ( .A0N(n1456), .A1N(n1453), .B0(n251), .Y(n1450) );
  OAI2BB1X1 U2672 ( .A0N(n1461), .A1N(n1459), .B0(n228), .Y(n1462) );
  OAI21XL U2673 ( .A0(n1459), .A1(work_cntr[10]), .B0(n1458), .Y(n1457) );
  OR2X1 U2674 ( .A(n132), .B(n1464), .Y(n1471) );
  OAI2BB1X1 U2675 ( .A0N(n1471), .A1N(n1468), .B0(n261), .Y(n1465) );
  OAI2BB1X1 U2676 ( .A0N(n1476), .A1N(n1474), .B0(n266), .Y(n1477) );
  OAI21XL U2677 ( .A0(n1474), .A1(work_cntr[8]), .B0(n140), .Y(n1472) );
  OAI21XL U2678 ( .A0(n1485), .A1(work_cntr[7]), .B0(n1488), .Y(n1486) );
  OA21XL U2679 ( .A0(n264), .A1(n1497), .B0(n1496), .Y(n1504) );
  OAI2BB1X1 U2680 ( .A0N(n1507), .A1N(n1501), .B0(n221), .Y(n1503) );
  OAI21XL U2681 ( .A0(n1501), .A1(work_cntr[5]), .B0(n1504), .Y(n1502) );
  OR2X1 U2682 ( .A(n1505), .B(n147), .Y(n1512) );
  OAI2BB1X1 U2683 ( .A0N(n1512), .A1N(n1510), .B0(n270), .Y(n1513) );
  OAI21XL U2684 ( .A0(n1510), .A1(work_cntr[4]), .B0(n1509), .Y(n1508) );
  OAI21XL U2685 ( .A0(n1520), .A1(N1827), .B0(n1522), .Y(n1521) );
  OAI22XL U2686 ( .A0(n1541), .A1(n1540), .B0(n1539), .B1(n1538), .Y(n1548) );
  OAI21XL U2687 ( .A0(N196), .A1(n1551), .B0(n1552), .Y(n1550) );
  NAND3BX1 U2688 ( .AN(write_cntr[12]), .B(n279), .C(n1558), .Y(n1561) );
  AOI2BB2X1 U2689 ( .B0(write_cntr[12]), .B1(n1560), .A0N(write_cntr[12]), 
        .A1N(n1560), .Y(n1565) );
  NAND3BX1 U2690 ( .AN(n1592), .B(write_cntr[7]), .C(n1588), .Y(n1577) );
  AOI2BB2X1 U2691 ( .B0(n1573), .B1(n1572), .A0N(n1573), .A1N(n1571), .Y(n1576) );
  NAND3BX1 U2692 ( .AN(n1628), .B(write_cntr[5]), .C(n1609), .Y(n1604) );
  AOI2BB2X1 U2693 ( .B0(n1600), .B1(n1599), .A0N(n1600), .A1N(n1599), .Y(n1613) );
  NAND3BX1 U2694 ( .AN(n1611), .B(n1613), .C(n1604), .Y(n1617) );
  AOI2BB2X1 U2695 ( .B0(n1603), .B1(n1602), .A0N(n1603), .A1N(n1601), .Y(n1615) );
  AOI2BB2X1 U2696 ( .B0(n1611), .B1(n1610), .A0N(n1611), .A1N(n1610), .Y(n1632) );
  AOI2BB2X1 U2697 ( .B0(n1609), .B1(n1608), .A0N(n1609), .A1N(n1608), .Y(n1634) );
  AOI2BB1X1 U2698 ( .A0N(n275), .A1N(n743), .B0(n1625), .Y(n1630) );
  OAI21XL U2699 ( .A0(write_cntr[4]), .A1(n1800), .B0(write_cntr[3]), .Y(n1626) );
  OAI221XL U2700 ( .A0(n1629), .A1(n1626), .B0(n1630), .B1(n1629), .C0(n1628), 
        .Y(n1627) );
  OAI31XL U2701 ( .A0(n1630), .A1(n1629), .A2(n1628), .B0(n1627), .Y(n1631) );
  OA21XL U2702 ( .A0(n1634), .A1(n1635), .B0(n1631), .Y(n1633) );
  AOI2BB1X1 U2703 ( .A0N(n1651), .A1N(n1650), .B0(n1659), .Y(n1654) );
  NAND3BX1 U2704 ( .AN(n1676), .B(n1664), .C(n1660), .Y(n1667) );
  AOI2BB2X1 U2705 ( .B0(n1666), .B1(n1665), .A0N(n1666), .A1N(n1664), .Y(n1668) );
  OAI21XL U2706 ( .A0(n1679), .A1(n1678), .B0(n1681), .Y(n1680) );
  AOI221XL U2707 ( .A0(n1698), .A1(n1692), .B0(n1699), .B1(n1692), .C0(n1702), 
        .Y(n1697) );
  AOI2BB2X1 U2708 ( .B0(n1694), .B1(n196), .A0N(n1694), .A1N(n196), .Y(n1696)
         );
  AOI2BB1X1 U2709 ( .A0N(n1697), .A1N(n1696), .B0(n1695), .Y(n1706) );
  OAI21XL U2710 ( .A0(n1704), .A1(n1700), .B0(n1702), .Y(n1701) );
  AO21X1 U2711 ( .A0(n1709), .A1(work_cntr[10]), .B0(n1705), .Y(n1716) );
  NAND3BX1 U2712 ( .AN(n1728), .B(n1720), .C(n1714), .Y(n1721) );
  OAI21XL U2713 ( .A0(n1720), .A1(n1719), .B0(n1718), .Y(n1722) );
  AO21X1 U2714 ( .A0(work_cntr[6]), .A1(n2446), .B0(n1730), .Y(n1735) );
  OAI2BB2XL U2715 ( .B0(n1738), .B1(n1737), .A0N(n1738), .A1N(n1737), .Y(n1740) );
  AO21X1 U2716 ( .A0(n1742), .A1(n1740), .B0(n1739), .Y(n1746) );
  AOI221XL U2717 ( .A0(n221), .A1(n2446), .B0(n1746), .B1(n2446), .C0(n1741), 
        .Y(n1743) );
  OAI21XL U2718 ( .A0(n1753), .A1(n1751), .B0(n1752), .Y(n1750) );
  OA22X1 U2719 ( .A0(n1767), .A1(n1766), .B0(n1765), .B1(n1764), .Y(n1768) );
  AOI2BB2X1 U2720 ( .B0(n1791), .B1(n1788), .A0N(n1773), .A1N(n1775), .Y(n1774) );
  ADDFXL U2721 ( .A(N1826), .B(n1777), .CI(n1776), .CO(n1778), .S(n1791) );
  AOI2BB2X1 U2722 ( .B0(n1779), .B1(n1778), .A0N(n1779), .A1N(n1778), .Y(n1792) );
  OAI31XL U2723 ( .A0(curr_photo_size[1]), .A1(n1784), .A2(n1787), .B0(n1796), 
        .Y(n1785) );
  AOI2BB2X1 U2724 ( .B0(n1813), .B1(n282), .A0N(n1813), .A1N(n282), .Y(n2782)
         );
  AOI2BB1X1 U2725 ( .A0N(write_addr[12]), .A1N(n1809), .B0(n1811), .Y(n2763)
         );
  AO21X1 U2726 ( .A0(n1815), .A1(n283), .B0(n1814), .Y(n2777) );
  AO21X1 U2727 ( .A0(n1818), .A1(n222), .B0(n1817), .Y(n2839) );
  AOI2BB2X1 U2728 ( .B0(n1835), .B1(n1834), .A0N(n1835), .A1N(n1834), .Y(n1842) );
  AOI2BB2X1 U2729 ( .B0(n1845), .B1(n1844), .A0N(n1845), .A1N(n1844), .Y(n1864) );
  AOI2BB2X1 U2730 ( .B0(n1850), .B1(n1849), .A0N(n1850), .A1N(n1849), .Y(n1865) );
  AOI2BB2X1 U2731 ( .B0(n1941), .B1(n1857), .A0N(n1856), .A1N(n1860), .Y(n1858) );
  AOI2BB2X1 U2732 ( .B0(n1859), .B1(n1858), .A0N(n1859), .A1N(n1858), .Y(n1885) );
  AOI2BB2X1 U2733 ( .B0(n131), .B1(n1876), .A0N(n131), .A1N(n1876), .Y(n1882)
         );
  OAI21XL U2734 ( .A0(n1929), .A1(n1880), .B0(n1877), .Y(n1878) );
  OAI22XL U2735 ( .A0(n1884), .A1(n1885), .B0(n1882), .B1(n1881), .Y(n1883) );
  OAI2BB1X1 U2736 ( .A0N(n1885), .A1N(n1884), .B0(n1883), .Y(n1891) );
  AOI2BB2X1 U2737 ( .B0(n1892), .B1(n174), .A0N(n1892), .A1N(n174), .Y(n1896)
         );
  AOI2BB2X1 U2738 ( .B0(n1928), .B1(n1896), .A0N(n1928), .A1N(n1896), .Y(n1893) );
  OAI22XL U2739 ( .A0(n2708), .A1(n1894), .B0(n1917), .B1(n1893), .Y(n1895) );
  AOI2BB2X1 U2740 ( .B0(n1900), .B1(n1899), .A0N(n1898), .A1N(n1906), .Y(n1911) );
  AOI2BB2X1 U2741 ( .B0(n1910), .B1(n1901), .A0N(n1910), .A1N(n1901), .Y(n1903) );
  AOI2BB2X1 U2742 ( .B0(n1924), .B1(n170), .A0N(n1924), .A1N(n170), .Y(n1914)
         );
  AOI2BB2X1 U2743 ( .B0(n1928), .B1(n1914), .A0N(n1928), .A1N(n1914), .Y(n1916) );
  AOI222XL U2744 ( .A0(n1928), .A1(n1924), .B0(n1928), .B1(n170), .C0(n1924), 
        .C1(n170), .Y(\intadd_3/CI ) );
  AOI2BB1X1 U2745 ( .A0N(n1926), .A1N(n2704), .B0(n1940), .Y(n1934) );
  ADDFXL U2746 ( .A(n1929), .B(n1928), .CI(n1927), .CO(n1930), .S(n1918) );
  AOI2BB1X1 U2747 ( .A0N(n1936), .A1N(next_cr_x[5]), .B0(n1943), .Y(n1939) );
  ADDFXL U2748 ( .A(n1936), .B(n1935), .CI(n1934), .CO(\intadd_3/B[2] ), .S(
        \intadd_3/A[1] ) );
  AOI2BB1X1 U2749 ( .A0N(n1941), .A1N(next_cr_x[6]), .B0(n2705), .Y(n1942) );
  ADDFXL U2750 ( .A(n1941), .B(n1940), .CI(n1939), .CO(\intadd_3/B[3] ), .S(
        \intadd_3/A[2] ) );
  ADDFXL U2751 ( .A(n2704), .B(n1943), .CI(n1942), .CO(\intadd_3/B[4] ), .S(
        \intadd_3/A[3] ) );
  AOI2BB2X1 U2752 ( .B0(n310), .B1(\intadd_3/SUM[4] ), .A0N(n2840), .A1N(n1944), .Y(n2852) );
  OAI21XL U2753 ( .A0(n2664), .A1(N1827), .B0(n2636), .Y(n1950) );
  OAI21XL U2754 ( .A0(n1972), .A1(n1971), .B0(n1970), .Y(n1967) );
  AOI2BB2X1 U2755 ( .B0(next_work_cntr[14]), .B1(n1969), .A0N(
        next_work_cntr[14]), .A1N(n1969), .Y(n1978) );
  OA21XL U2756 ( .A0(n1972), .A1(n1971), .B0(n1970), .Y(n1975) );
  OAI21XL U2757 ( .A0(n1975), .A1(n1974), .B0(n1973), .Y(n1977) );
  AOI2BB2X1 U2758 ( .B0(n1982), .B1(n1981), .A0N(n1982), .A1N(n1981), .Y(n1984) );
  AO21X1 U2759 ( .A0(n1992), .A1(n1991), .B0(n1990), .Y(n1994) );
  AOI2BB2X1 U2760 ( .B0(n2001), .B1(n169), .A0N(n2001), .A1N(n169), .Y(n2002)
         );
  OAI31XL U2761 ( .A0(n2003), .A1(n2008), .A2(n168), .B0(n2002), .Y(n2005) );
  AOI2BB2X1 U2762 ( .B0(next_work_cntr[10]), .B1(n2009), .A0N(
        next_work_cntr[10]), .A1N(n2009), .Y(n2021) );
  OAI21XL U2763 ( .A0(n2033), .A1(n2032), .B0(n2017), .Y(n2024) );
  AOI2BB2X1 U2764 ( .B0(n2031), .B1(n2030), .A0N(n2031), .A1N(n2030), .Y(n2038) );
  AOI2BB2X1 U2765 ( .B0(n2045), .B1(n2057), .A0N(n2045), .A1N(n2057), .Y(n2058) );
  OAI21XL U2766 ( .A0(n2049), .A1(n2048), .B0(n2047), .Y(n2050) );
  AOI2BB2X1 U2767 ( .B0(n2065), .B1(n2064), .A0N(n2065), .A1N(n2064), .Y(n2067) );
  OAI21XL U2768 ( .A0(n2099), .A1(n2102), .B0(n2091), .Y(n2088) );
  OAI22XL U2769 ( .A0(n2100), .A1(n2088), .B0(n2099), .B1(n2091), .Y(n2105) );
  AOI221XL U2770 ( .A0(n2099), .A1(n2093), .B0(n2102), .B1(n2093), .C0(n2092), 
        .Y(n2094) );
  OAI21XL U2771 ( .A0(n2098), .A1(n2094), .B0(n2096), .Y(n2095) );
  OAI21XL U2772 ( .A0(n2100), .A1(n2099), .B0(n2103), .Y(n2101) );
  OAI21XL U2773 ( .A0(n2103), .A1(n2102), .B0(n2101), .Y(n2104) );
  NAND3BX1 U2774 ( .AN(n2112), .B(n2118), .C(n2128), .Y(n2119) );
  AO21X1 U2775 ( .A0(next_work_cntr[14]), .A1(n2117), .B0(n130), .Y(n2157) );
  AOI2BB2X1 U2776 ( .B0(next_work_cntr[15]), .B1(n130), .A0N(
        next_work_cntr[15]), .A1N(n130), .Y(n2159) );
  AND4X1 U2777 ( .A(n2153), .B(n2137), .C(n2191), .D(n2189), .Y(n2126) );
  NAND3BX1 U2778 ( .AN(n2151), .B(n2172), .C(n2126), .Y(n2138) );
  OR2X1 U2779 ( .A(n2140), .B(n2138), .Y(n2141) );
  AO21X1 U2780 ( .A0(n2135), .A1(n2134), .B0(n2133), .Y(n2160) );
  AOI2BB2X1 U2781 ( .B0(n2140), .B1(n2139), .A0N(n2140), .A1N(n2139), .Y(n2142) );
  AOI2BB2X1 U2782 ( .B0(n2155), .B1(n2149), .A0N(n2155), .A1N(n2149), .Y(n2177) );
  NOR4X1 U2783 ( .A(n2178), .B(next_work_cntr[7]), .C(n2151), .D(n2150), .Y(
        n2179) );
  OAI21XL U2784 ( .A0(n2158), .A1(n2176), .B0(n2157), .Y(n2156) );
  NAND3BX1 U2785 ( .AN(n2159), .B(n2179), .C(n2188), .Y(n2196) );
  OAI21XL U2786 ( .A0(n2173), .A1(n2175), .B0(n2172), .Y(n2171) );
  OAI22XL U2787 ( .A0(n2209), .A1(n2207), .B0(n2193), .B1(n2192), .Y(n2194) );
  OR2X1 U2788 ( .A(n2214), .B(n2215), .Y(n2206) );
  AOI2BB2X1 U2789 ( .B0(n2209), .B1(n2208), .A0N(n2209), .A1N(n2208), .Y(n2252) );
  OR2X1 U2790 ( .A(n2211), .B(n2210), .Y(n2213) );
  AOI2BB2X1 U2791 ( .B0(n2215), .B1(n2214), .A0N(n2215), .A1N(n2214), .Y(n2248) );
  OAI21XL U2792 ( .A0(n2241), .A1(n2242), .B0(n2243), .Y(n2240) );
  AOI2BB2X1 U2793 ( .B0(n2245), .B1(n2244), .A0N(n2245), .A1N(n2244), .Y(n2269) );
  NAND3BX1 U2794 ( .AN(n2275), .B(n2266), .C(n210), .Y(n2270) );
  AOI2BB1X1 U2795 ( .A0N(next_work_cntr[3]), .A1N(n2270), .B0(n2304), .Y(n2302) );
  OAI21XL U2796 ( .A0(n2278), .A1(n2295), .B0(n2277), .Y(n2276) );
  OAI21XL U2797 ( .A0(n2286), .A1(n2285), .B0(n2309), .Y(n2284) );
  OAI21XL U2798 ( .A0(n211), .A1(n2297), .B0(n2298), .Y(n2296) );
  OAI31XL U2799 ( .A0(n211), .A1(n2298), .A2(n2297), .B0(n2296), .Y(n2299) );
  OAI21XL U2800 ( .A0(n2310), .A1(n2309), .B0(n2314), .Y(n2311) );
  AOI2BB2X1 U2801 ( .B0(n2312), .B1(n2331), .A0N(n2312), .A1N(n2331), .Y(n2328) );
  AOI2BB2X1 U2802 ( .B0(n2319), .B1(n2318), .A0N(n2319), .A1N(n2318), .Y(n2322) );
  AOI2BB2X1 U2803 ( .B0(n2322), .B1(n2321), .A0N(n2322), .A1N(n2321), .Y(n2346) );
  AOI2BB2X1 U2804 ( .B0(next_work_cntr[1]), .B1(n2327), .A0N(next_work_cntr[1]), .A1N(n2327), .Y(n2353) );
  AOI2BB2X1 U2805 ( .B0(n2334), .B1(n2364), .A0N(n2334), .A1N(n2364), .Y(n2357) );
  AOI2BB2X1 U2806 ( .B0(n2336), .B1(n2335), .A0N(n2336), .A1N(n2335), .Y(n2363) );
  OAI21XL U2807 ( .A0(n2344), .A1(n2346), .B0(n2347), .Y(n2345) );
  NAND4BBXL U2808 ( .AN(n2357), .BN(n2356), .C(n2355), .D(n2354), .Y(n2360) );
  OAI31XL U2809 ( .A0(n2366), .A1(n2365), .A2(n2364), .B0(n2363), .Y(n2367) );
  AOI222XL U2810 ( .A0(n2804), .A1(n2377), .B0(n2804), .B1(n2376), .C0(n2377), 
        .C1(n2375), .Y(n2678) );
  AO21X1 U2811 ( .A0(n2394), .A1(work_cntr[17]), .B0(n2387), .Y(n2388) );
  AO21X1 U2812 ( .A0(n2389), .A1(n2390), .B0(n2391), .Y(n2402) );
  OR2X1 U2813 ( .A(n2389), .B(n2390), .Y(n2392) );
  AOI222XL U2814 ( .A0(n2399), .A1(n2400), .B0(n2399), .B1(n2396), .C0(n2400), 
        .C1(work_cntr[16]), .Y(n2397) );
  AOI2BB2X1 U2815 ( .B0(n2398), .B1(n2397), .A0N(n2398), .A1N(n2401), .Y(n2405) );
  OAI21XL U2816 ( .A0(work_cntr[14]), .A1(n2412), .B0(n2420), .Y(n2408) );
  NOR3BXL U2817 ( .AN(n2421), .B(n2418), .C(n2420), .Y(n2411) );
  OAI2BB1X1 U2818 ( .A0N(n2413), .A1N(n2425), .B0(n2430), .Y(n2429) );
  OAI2BB1X1 U2819 ( .A0N(n2416), .A1N(work_cntr[12]), .B0(n2415), .Y(n2435) );
  OAI21XL U2820 ( .A0(n2418), .A1(n2420), .B0(n2421), .Y(n2419) );
  AO21X1 U2821 ( .A0(n2423), .A1(n2428), .B0(n2422), .Y(n2424) );
  AO21X1 U2822 ( .A0(n217), .A1(n2439), .B0(n2436), .Y(n2427) );
  AOI2BB2X1 U2823 ( .B0(n2429), .B1(n2428), .A0N(n2429), .A1N(n2427), .Y(n2437) );
  AO21X1 U2824 ( .A0(n251), .A1(n2444), .B0(n2437), .Y(n2438) );
  AOI2BB2X1 U2825 ( .B0(n2440), .B1(n2439), .A0N(n2440), .A1N(n2438), .Y(n2451) );
  OAI21XL U2826 ( .A0(work_cntr[10]), .A1(n2453), .B0(n2445), .Y(n2442) );
  AOI2BB2X1 U2827 ( .B0(n2443), .B1(n2444), .A0N(n2443), .A1N(n2442), .Y(n2452) );
  OR2X1 U2828 ( .A(n2445), .B(n2444), .Y(n2449) );
  AOI2BB1X1 U2829 ( .A0N(n2448), .A1N(n266), .B0(n2447), .Y(n2455) );
  AOI2BB2X1 U2830 ( .B0(n268), .B1(n2464), .A0N(n268), .A1N(n2464), .Y(n2458)
         );
  AO21X1 U2831 ( .A0(n266), .A1(n2468), .B0(n2463), .Y(n2454) );
  AOI2BB2X1 U2832 ( .B0(n2456), .B1(n2455), .A0N(n2456), .A1N(n2454), .Y(n2466) );
  OA21XL U2833 ( .A0(n2466), .A1(n2458), .B0(n2474), .Y(n2473) );
  OA21XL U2834 ( .A0(n2463), .A1(n2462), .B0(n2461), .Y(n2469) );
  AO21X1 U2835 ( .A0(n268), .A1(n2471), .B0(n2466), .Y(n2467) );
  OAI21XL U2836 ( .A0(work_cntr[6]), .A1(n164), .B0(n2470), .Y(n2472) );
  AOI2BB2X1 U2837 ( .B0(n2473), .B1(n2472), .A0N(n2473), .A1N(n2471), .Y(n2483) );
  OA21XL U2838 ( .A0(n2483), .A1(n164), .B0(n2478), .Y(n2490) );
  OAI21XL U2839 ( .A0(n2484), .A1(n221), .B0(n2478), .Y(n2488) );
  OAI21XL U2840 ( .A0(work_cntr[5]), .A1(n2484), .B0(n2483), .Y(n2485) );
  OAI21XL U2841 ( .A0(work_cntr[4]), .A1(n2503), .B0(n2494), .Y(n2489) );
  AOI2BB2X1 U2842 ( .B0(n2490), .B1(n2495), .A0N(n2490), .A1N(n2489), .Y(n2493) );
  AOI2BB2X1 U2843 ( .B0(n2495), .B1(n2494), .A0N(n2495), .A1N(n2494), .Y(n2502) );
  OAI21XL U2844 ( .A0(n2498), .A1(n2503), .B0(n2502), .Y(n2501) );
  AOI2BB2X1 U2845 ( .B0(N1826), .B1(n2507), .A0N(N1826), .A1N(n2507), .Y(n2509) );
  AO21X1 U2846 ( .A0(n2511), .A1(N1825), .B0(N196), .Y(n2508) );
  OAI21XL U2847 ( .A0(n2511), .A1(N1825), .B0(n2510), .Y(n2512) );
  NAND3BX1 U2848 ( .AN(n2522), .B(n2521), .C(n2520), .Y(n2528) );
  OAI2BB1X1 U2849 ( .A0N(n2524), .A1N(n2528), .B0(n2526), .Y(n2530) );
  OAI21XL U2850 ( .A0(n2528), .A1(n2527), .B0(n2531), .Y(n2529) );
  OR2X1 U2851 ( .A(n2532), .B(n2537), .Y(n2541) );
  OAI2BB1X1 U2852 ( .A0N(n2541), .A1N(n2536), .B0(n2539), .Y(n2538) );
  OAI2BB1X1 U2853 ( .A0N(n2543), .A1N(n2546), .B0(n2545), .Y(n2547) );
  OR2X1 U2854 ( .A(n2549), .B(n2554), .Y(n2558) );
  OAI2BB1X1 U2855 ( .A0N(n2558), .A1N(n2553), .B0(n2556), .Y(n2555) );
  OAI31XL U2856 ( .A0(n2553), .A1(n2552), .A2(n2551), .B0(n2550), .Y(n2559) );
  OAI2BB1X1 U2857 ( .A0N(n2560), .A1N(n2564), .B0(n2562), .Y(n2566) );
  OAI21XL U2858 ( .A0(n2564), .A1(n2563), .B0(n2567), .Y(n2565) );
  OR2X1 U2859 ( .A(n2573), .B(n2568), .Y(n2577) );
  OAI2BB1X1 U2860 ( .A0N(n2577), .A1N(n2572), .B0(n2575), .Y(n2574) );
  OA21XL U2861 ( .A0(n2575), .A1(n2576), .B0(n2574), .Y(n2586) );
  OAI2BB1X1 U2862 ( .A0N(n2579), .A1N(n2583), .B0(n2581), .Y(n2585) );
  OAI21XL U2863 ( .A0(n2583), .A1(n2582), .B0(n2586), .Y(n2584) );
  OR2X1 U2864 ( .A(n143), .B(n2587), .Y(n2596) );
  OAI2BB1X1 U2865 ( .A0N(n2596), .A1N(n2591), .B0(n2594), .Y(n2593) );
  OAI2BB1X1 U2866 ( .A0N(n2598), .A1N(n2602), .B0(n2600), .Y(n2604) );
  OAI21XL U2867 ( .A0(n2602), .A1(n2601), .B0(n2605), .Y(n2603) );
  OR2X1 U2868 ( .A(n2611), .B(n2606), .Y(n2615) );
  OAI2BB1X1 U2869 ( .A0N(n2615), .A1N(n2610), .B0(n2613), .Y(n2612) );
  OA21XL U2870 ( .A0(n2613), .A1(n2614), .B0(n2612), .Y(n2624) );
  OAI2BB1X1 U2871 ( .A0N(n2617), .A1N(n2621), .B0(n2619), .Y(n2623) );
  OAI21XL U2872 ( .A0(n2621), .A1(n2620), .B0(n2624), .Y(n2622) );
  OR2X1 U2873 ( .A(n145), .B(n2625), .Y(n2631) );
  OAI2BB1X1 U2874 ( .A0N(n2631), .A1N(n2629), .B0(n2634), .Y(n2632) );
  OA21XL U2875 ( .A0(n2634), .A1(n2633), .B0(n2632), .Y(n2641) );
  OAI2BB1X1 U2876 ( .A0N(n2645), .A1N(n2638), .B0(n2636), .Y(n2640) );
  OAI21XL U2877 ( .A0(n2638), .A1(n2637), .B0(n2641), .Y(n2639) );
  OR2X1 U2878 ( .A(n144), .B(n2643), .Y(n2651) );
  OAI2BB1X1 U2879 ( .A0N(n2651), .A1N(n2649), .B0(n2654), .Y(n2652) );
  OAI21XL U2880 ( .A0(n2649), .A1(n2646), .B0(n2648), .Y(n2647) );
  OA21XL U2881 ( .A0(n2672), .A1(n2668), .B0(n2666), .Y(n2670) );
  AOI2BB2X1 U2882 ( .B0(n2672), .B1(n2667), .A0N(n2672), .A1N(n2667), .Y(n2675) );
  OAI2BB1X1 U2883 ( .A0N(n2668), .A1N(n2669), .B0(n2667), .Y(n2671) );
  OAI2BB2XL U2884 ( .B0(n2670), .B1(n2669), .A0N(n284), .A1N(n2671), .Y(n2674)
         );
  AOI2BB1X1 U2885 ( .A0N(N196), .A1N(n2672), .B0(n2671), .Y(n2673) );
  AO21X1 U2886 ( .A0(n2689), .A1(n302), .B0(n2699), .Y(n2691) );
  OAI2BB1X1 U2887 ( .A0N(n2694), .A1N(cr_read_cntr[5]), .B0(n2693), .Y(n449)
         );
  AOI2BB1X1 U2888 ( .A0N(cr_read_cntr[6]), .A1N(n2697), .B0(n2698), .Y(n448)
         );
  OA21XL U2889 ( .A0(cr_read_cntr[7]), .A1(n2700), .B0(n2701), .Y(n447) );
  ADDFXL U2890 ( .A(next_cr_x[5]), .B(n2705), .CI(n2704), .CO(\intadd_3/B[5] ), 
        .S(\intadd_3/A[4] ) );
  OAI2BB2XL U2891 ( .B0(n2771), .B1(n235), .A0N(n310), .A1N(\intadd_3/SUM[5] ), 
        .Y(n2706) );
  ADDFXL U2892 ( .A(n230), .B(next_cr_x[6]), .CI(n2712), .CO(\intadd_3/B[7] ), 
        .S(\intadd_3/B[6] ) );
  NAND3BX1 U2893 ( .AN(n2734), .B(n2730), .C(n2731), .Y(n2729) );
  AOI2BB2X1 U2894 ( .B0(n2738), .B1(n2737), .A0N(n2738), .A1N(n2736), .Y(n2745) );
  AOI2BB2X1 U2895 ( .B0(n2745), .B1(n2744), .A0N(n2745), .A1N(n2743), .Y(n2750) );
  AOI2BB2X1 U2896 ( .B0(n2753), .B1(n2752), .A0N(n2753), .A1N(n2751), .Y(n2760) );
  AOI2BB2X1 U2897 ( .B0(n2758), .B1(n2754), .A0N(n2758), .A1N(n2759), .Y(
        \intadd_3/B[8] ) );
  AO21X1 U2898 ( .A0(n310), .A1(\intadd_3/SUM[8] ), .B0(n2757), .Y(n2858) );
  AO22X1 U2899 ( .A0(n2761), .A1(n2760), .B0(n2759), .B1(n2758), .Y(
        \intadd_3/A[9] ) );
  OAI21XL U2900 ( .A0(n2763), .A1(n2762), .B0(n2765), .Y(n2764) );
  AO21X1 U2901 ( .A0(n246), .A1(n310), .B0(n2767), .Y(n2828) );
  AOI2BB2X1 U2902 ( .B0(n2770), .B1(n2775), .A0N(n2770), .A1N(n2775), .Y(n2772) );
  NAND3BX1 U2903 ( .AN(n2775), .B(n2774), .C(n2773), .Y(n2776) );
  AOI2BB2X1 U2904 ( .B0(curr_photo[1]), .B1(photo_num[1]), .A0N(curr_photo[1]), 
        .A1N(photo_num[1]), .Y(n2788) );
  AOI2BB2X1 U2905 ( .B0(curr_photo[0]), .B1(photo_num[0]), .A0N(curr_photo[0]), 
        .A1N(photo_num[0]), .Y(n2787) );
  OAI21XL U2906 ( .A0(n2804), .A1(n2798), .B0(n285), .Y(n2799) );
  OAI21XL U2907 ( .A0(n2804), .A1(write_addr[8]), .B0(n2809), .Y(n2805) );
  OR2X1 U2908 ( .A(n2820), .B(n2853), .Y(n2823) );
endmodule


module DPA ( clk, reset, IM_A, IM_Q, IM_D, IM_WEN, CR_A, CR_Q );
  output [19:0] IM_A;
  input [23:0] IM_Q;
  output [23:0] IM_D;
  output [8:0] CR_A;
  input [12:0] CR_Q;
  input clk, reset;
  output IM_WEN;
  wire   n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         im_d_w_19, im_d_w_18, im_d_w_9, im_d_w_8, en_si, en_init_time,
         en_photo_num, en_curr_photo_size, en_so, si_sel, init_time_mux_sel,
         \sftr_n[0] , \data_path/si_w[0] , \data_path/si_w[1] ,
         \data_path/si_w[2] , \data_path/si_w[3] , \data_path/si_w[4] ,
         \data_path/si_w[5] , \data_path/si_w[6] , \data_path/si_w[7] ,
         \data_path/si_w[8] , \data_path/si_w[9] , \data_path/si_w[10] ,
         \data_path/si_w[11] , \data_path/si_w[12] , \data_path/si_w[13] ,
         \data_path/si_w[14] , \data_path/si_w[15] , \data_path/si_w[16] ,
         \data_path/si_w[17] , \data_path/si_w[18] , \data_path/si_w[19] ,
         \data_path/si_w[20] , \data_path/si_w[21] , \data_path/si_w[22] ,
         \data_path/si_w[23] , n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n141, n144, n145, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, \intadd_0/CI , \intadd_0/SUM[6] ,
         \intadd_0/SUM[5] , \intadd_0/SUM[4] , \intadd_0/SUM[3] ,
         \intadd_0/SUM[2] , \intadd_0/SUM[1] , \intadd_0/SUM[0] ,
         \intadd_0/n7 , \intadd_0/n6 , \intadd_0/n5 , \intadd_0/n4 ,
         \intadd_0/n3 , \intadd_0/n2 , \intadd_0/n1 , \intadd_1/CI ,
         \intadd_1/SUM[6] , \intadd_1/SUM[5] , \intadd_1/SUM[4] ,
         \intadd_1/SUM[3] , \intadd_1/SUM[2] , \intadd_1/SUM[1] ,
         \intadd_1/SUM[0] , \intadd_1/n7 , \intadd_1/n6 , \intadd_1/n5 ,
         \intadd_1/n4 , \intadd_1/n3 , \intadd_1/n2 , \intadd_1/n1 ,
         \intadd_2/CI , \intadd_2/SUM[6] , \intadd_2/SUM[5] ,
         \intadd_2/SUM[4] , \intadd_2/SUM[3] , \intadd_2/SUM[2] ,
         \intadd_2/SUM[1] , \intadd_2/SUM[0] , \intadd_2/n7 , \intadd_2/n6 ,
         \intadd_2/n5 , \intadd_2/n4 , \intadd_2/n3 , \intadd_2/n2 ,
         \intadd_2/n1 , n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n442, n444, n446, n448, n450, n452, n454, n456, n458, n460, n462,
         n464, n465, n466, n467, n468, n469, n470, n471, n473, n475, n477,
         n480, n482, n484, n486, n488, n490, n492, n494, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n754;
  wire   [29:28] im_d_w;
  wire   [23:0] curr_time;
  wire   [19:0] fb_addr;
  wire   [1:0] photo_num;
  wire   [19:0] curr_photo_addr;
  wire   [1:0] curr_photo_size;
  wire   [1:0] so_mux_sel;
  wire   [3:0] expand_sel;

  CONT ctrl_logic ( .clk(clk), .reset(reset), .im_wen_n(IM_WEN), .cr_a(CR_A), 
        .curr_time({curr_time[23:3], n470, curr_time[1:0]}), .fb_addr(fb_addr), 
        .photo_num(photo_num), .curr_photo_addr(curr_photo_addr), 
        .curr_photo_size(curr_photo_size), .en_si(en_si), .en_init_time(
        en_init_time), .en_fb_addr(n468), .en_photo_num(en_photo_num), 
        .en_curr_photo_addr(n469), .en_curr_photo_size(en_curr_photo_size), 
        .en_so(en_so), .si_sel(si_sel), .init_time_mux_sel(init_time_mux_sel), 
        .so_mux_sel(so_mux_sel), .expand_sel(expand_sel), .\im_a[19]_BAR (n755), .\im_a[18]_BAR (n756), .\im_a[17]_BAR (n757), .\im_a[16]_BAR (n758), 
        .\im_a[15]_BAR (n759), .\im_a[14]_BAR (n760), .\im_a[13]_BAR (n761), 
        .\im_a[12]_BAR (n762), .\im_a[11]_BAR (n763), .\im_a[10]_BAR (n764), 
        .\im_a[9]_BAR (n765), .\im_a[8]_BAR (n766), .\im_a[7]_BAR (n767), 
        .\im_a[6]_BAR (n768), .\im_a[5]_BAR (n769), .\im_a[4]_BAR (n770), 
        .\im_a[3]_BAR (n771), .\im_a[2]_BAR (n772), .\im_a[1]_BAR (n773), 
        .\im_a[0]_BAR (n774), .\sftr_n[0]_BAR (\sftr_n[0] ) );
  ADDFXL \intadd_0/U3  ( .A(n776), .B(\data_path/si_w[22] ), .CI(\intadd_0/n3 ), .CO(\intadd_0/n2 ), .S(\intadd_0/SUM[5] ) );
  ADDFXL \intadd_1/U3  ( .A(IM_D[14]), .B(\data_path/si_w[14] ), .CI(
        \intadd_1/n3 ), .CO(\intadd_1/n2 ), .S(\intadd_1/SUM[5] ) );
  ADDFXL \intadd_2/U3  ( .A(IM_D[6]), .B(\data_path/si_w[6] ), .CI(
        \intadd_2/n3 ), .CO(\intadd_2/n2 ), .S(\intadd_2/SUM[5] ) );
  DFFSX1 \data_path/si_reg/q_reg[2]  ( .D(n314), .CK(clk), .SN(n542), .Q(n510), 
        .QN(\data_path/si_w[2] ) );
  DFFSX1 \data_path/si_reg/q_reg[4]  ( .D(n313), .CK(clk), .SN(n542), .Q(n509), 
        .QN(\data_path/si_w[4] ) );
  DFFSX1 \data_path/si_reg/q_reg[1]  ( .D(n315), .CK(clk), .SN(n22), .Q(n504), 
        .QN(\data_path/si_w[1] ) );
  DFFSX1 \data_path/si_reg/q_reg[8]  ( .D(n312), .CK(clk), .SN(n542), .Q(n500), 
        .QN(\data_path/si_w[8] ) );
  DFFSX1 \data_path/init_time_reg/q_reg[1]  ( .D(n145), .CK(clk), .SN(n542), 
        .Q(n649), .QN(curr_time[1]) );
  ADDFXL \intadd_2/U7  ( .A(IM_D[2]), .B(\data_path/si_w[2] ), .CI(
        \intadd_2/n7 ), .CO(\intadd_2/n6 ), .S(\intadd_2/SUM[1] ) );
  ADDFXL \intadd_2/U2  ( .A(IM_D[7]), .B(\data_path/si_w[7] ), .CI(
        \intadd_2/n2 ), .CO(\intadd_2/n1 ), .S(\intadd_2/SUM[6] ) );
  ADDFXL \intadd_1/U7  ( .A(n785), .B(\data_path/si_w[10] ), .CI(\intadd_1/n7 ), .CO(\intadd_1/n6 ), .S(\intadd_1/SUM[1] ) );
  ADDFXL \intadd_1/U2  ( .A(IM_D[15]), .B(\data_path/si_w[15] ), .CI(
        \intadd_1/n2 ), .CO(\intadd_1/n1 ), .S(\intadd_1/SUM[6] ) );
  ADDFXL \intadd_0/U7  ( .A(IM_D[18]), .B(\data_path/si_w[18] ), .CI(
        \intadd_0/n7 ), .CO(\intadd_0/n6 ), .S(\intadd_0/SUM[1] ) );
  ADDFXL \intadd_0/U2  ( .A(n775), .B(\data_path/si_w[23] ), .CI(\intadd_0/n2 ), .CO(\intadd_0/n1 ), .S(\intadd_0/SUM[6] ) );
  ADDFXL \intadd_1/U8  ( .A(n786), .B(\data_path/si_w[9] ), .CI(\intadd_1/CI ), 
        .CO(\intadd_1/n7 ), .S(\intadd_1/SUM[0] ) );
  ADDFXL \intadd_0/U8  ( .A(n781), .B(\data_path/si_w[17] ), .CI(\intadd_0/CI ), .CO(\intadd_0/n7 ), .S(\intadd_0/SUM[0] ) );
  ADDFXL \intadd_2/U8  ( .A(IM_D[1]), .B(\data_path/si_w[1] ), .CI(
        \intadd_2/CI ), .CO(\intadd_2/n7 ), .S(\intadd_2/SUM[0] ) );
  ADDFXL \intadd_2/U6  ( .A(IM_D[3]), .B(\data_path/si_w[3] ), .CI(
        \intadd_2/n6 ), .CO(\intadd_2/n5 ), .S(\intadd_2/SUM[2] ) );
  ADDFXL \intadd_2/U5  ( .A(IM_D[4]), .B(\data_path/si_w[4] ), .CI(
        \intadd_2/n5 ), .CO(\intadd_2/n4 ), .S(\intadd_2/SUM[3] ) );
  ADDFXL \intadd_2/U4  ( .A(IM_D[5]), .B(\data_path/si_w[5] ), .CI(
        \intadd_2/n4 ), .CO(\intadd_2/n3 ), .S(\intadd_2/SUM[4] ) );
  ADDFXL \intadd_1/U6  ( .A(n784), .B(\data_path/si_w[11] ), .CI(\intadd_1/n6 ), .CO(\intadd_1/n5 ), .S(\intadd_1/SUM[2] ) );
  ADDFXL \intadd_1/U5  ( .A(n783), .B(\data_path/si_w[12] ), .CI(\intadd_1/n5 ), .CO(\intadd_1/n4 ), .S(\intadd_1/SUM[3] ) );
  ADDFXL \intadd_1/U4  ( .A(IM_D[13]), .B(\data_path/si_w[13] ), .CI(
        \intadd_1/n4 ), .CO(\intadd_1/n3 ), .S(\intadd_1/SUM[4] ) );
  ADDFXL \intadd_0/U6  ( .A(n779), .B(\data_path/si_w[19] ), .CI(\intadd_0/n6 ), .CO(\intadd_0/n5 ), .S(\intadd_0/SUM[2] ) );
  ADDFXL \intadd_0/U5  ( .A(n778), .B(\data_path/si_w[20] ), .CI(\intadd_0/n5 ), .CO(\intadd_0/n4 ), .S(\intadd_0/SUM[3] ) );
  ADDFXL \intadd_0/U4  ( .A(n777), .B(\data_path/si_w[21] ), .CI(\intadd_0/n4 ), .CO(\intadd_0/n3 ), .S(\intadd_0/SUM[4] ) );
  DFFSX2 \data_path/init_time_reg/q_reg[4]  ( .D(n141), .CK(clk), .SN(n542), 
        .QN(curr_time[4]) );
  DFFSX2 \data_path/init_time_reg/q_reg[2]  ( .D(n144), .CK(clk), .SN(n22), 
        .QN(n470) );
  DFFRX2 \data_path/si_reg/q_reg[16]  ( .D(n418), .CK(clk), .RN(n22), .Q(
        \data_path/si_w[16] ) );
  DFFRX2 \data_path/init_time_reg/q_reg[15]  ( .D(n324), .CK(clk), .RN(n22), 
        .Q(curr_time[15]) );
  DFFRX2 \data_path/init_time_reg/q_reg[14]  ( .D(n325), .CK(clk), .RN(n22), 
        .Q(curr_time[14]) );
  DFFRX2 \data_path/init_time_reg/q_reg[7]  ( .D(n332), .CK(clk), .RN(n22), 
        .Q(curr_time[7]) );
  DFFRX2 \data_path/init_time_reg/q_reg[6]  ( .D(n333), .CK(clk), .RN(n22), 
        .Q(curr_time[6]) );
  DFFRX2 \data_path/init_time_reg/q_reg[17]  ( .D(n322), .CK(clk), .RN(n22), 
        .Q(curr_time[17]), .QN(n679) );
  DFFRX2 \data_path/si_reg/q_reg[0]  ( .D(n417), .CK(clk), .RN(n22), .Q(
        \data_path/si_w[0] ), .QN(n498) );
  DFFRX2 \data_path/curr_photo_size_reg/q_reg[0]  ( .D(n368), .CK(clk), .RN(
        n22), .Q(curr_photo_size[0]), .QN(n514) );
  DFFRX2 \data_path/init_time_reg/q_reg[9]  ( .D(n330), .CK(clk), .RN(n22), 
        .Q(curr_time[9]), .QN(n529) );
  DFFRX2 \data_path/init_time_reg/q_reg[12]  ( .D(n327), .CK(clk), .RN(n22), 
        .Q(curr_time[12]), .QN(n518) );
  DFFRX2 \data_path/init_time_reg/q_reg[10]  ( .D(n329), .CK(clk), .RN(n22), 
        .Q(curr_time[10]), .QN(n505) );
  DFFRX1 \data_path/si_reg/q_reg[23]  ( .D(n369), .CK(clk), .RN(n22), .Q(
        \data_path/si_w[23] ), .QN(n513) );
  DFFRX1 \data_path/si_reg/q_reg[22]  ( .D(n370), .CK(clk), .RN(n22), .Q(
        \data_path/si_w[22] ), .QN(n512) );
  DFFRX1 \data_path/si_reg/q_reg[21]  ( .D(n371), .CK(clk), .RN(n22), .Q(
        \data_path/si_w[21] ), .QN(n511) );
  DFFRX1 \data_path/si_reg/q_reg[20]  ( .D(n372), .CK(clk), .RN(n542), .Q(
        \data_path/si_w[20] ), .QN(n532) );
  DFFRX1 \data_path/si_reg/q_reg[19]  ( .D(n375), .CK(clk), .RN(n542), .Q(
        \data_path/si_w[19] ), .QN(n526) );
  DFFRX1 \data_path/si_reg/q_reg[18]  ( .D(n378), .CK(clk), .RN(n467), .Q(
        \data_path/si_w[18] ), .QN(n524) );
  DFFRX1 \data_path/si_reg/q_reg[17]  ( .D(n381), .CK(clk), .RN(n467), .Q(
        \data_path/si_w[17] ), .QN(n525) );
  DFFRX1 \data_path/si_reg/q_reg[15]  ( .D(n384), .CK(clk), .RN(n467), .Q(
        \data_path/si_w[15] ), .QN(n523) );
  DFFRX1 \data_path/si_reg/q_reg[14]  ( .D(n387), .CK(clk), .RN(n467), .Q(
        \data_path/si_w[14] ), .QN(n527) );
  DFFRX1 \data_path/si_reg/q_reg[13]  ( .D(n390), .CK(clk), .RN(n467), .Q(
        \data_path/si_w[13] ), .QN(n507) );
  DFFRX1 \data_path/si_reg/q_reg[12]  ( .D(n393), .CK(clk), .RN(n22), .Q(
        \data_path/si_w[12] ), .QN(n520) );
  DFFRX1 \data_path/si_reg/q_reg[11]  ( .D(n396), .CK(clk), .RN(n22), .Q(
        \data_path/si_w[11] ), .QN(n501) );
  DFFRX1 \data_path/si_reg/q_reg[10]  ( .D(n399), .CK(clk), .RN(n542), .Q(
        \data_path/si_w[10] ), .QN(n499) );
  DFFRX1 \data_path/si_reg/q_reg[9]  ( .D(n402), .CK(clk), .RN(n542), .Q(
        \data_path/si_w[9] ), .QN(n521) );
  DFFRX1 \data_path/si_reg/q_reg[7]  ( .D(n405), .CK(clk), .RN(n542), .Q(
        \data_path/si_w[7] ), .QN(n517) );
  DFFRX1 \data_path/si_reg/q_reg[6]  ( .D(n408), .CK(clk), .RN(n467), .Q(
        \data_path/si_w[6] ), .QN(n522) );
  DFFRX1 \data_path/si_reg/q_reg[5]  ( .D(n411), .CK(clk), .RN(n467), .Q(
        \data_path/si_w[5] ), .QN(n508) );
  DFFRX1 \data_path/si_reg/q_reg[3]  ( .D(n414), .CK(clk), .RN(n467), .Q(
        \data_path/si_w[3] ), .QN(n516) );
  DFFRX1 \data_path/photo_num_reg/q_reg[1]  ( .D(n21), .CK(clk), .RN(n542), 
        .Q(photo_num[1]), .QN(n10) );
  DFFRX1 \data_path/curr_photo_size_reg/q_reg[1]  ( .D(n23), .CK(clk), .RN(n22), .Q(curr_photo_size[1]), .QN(n530) );
  DFFRX1 \data_path/init_time_reg/q_reg[16]  ( .D(n323), .CK(clk), .RN(n22), 
        .Q(curr_time[16]), .QN(n506) );
  DFFRX1 \data_path/init_time_reg/q_reg[19]  ( .D(n320), .CK(clk), .RN(n542), 
        .Q(curr_time[19]), .QN(n535) );
  DFFRX1 \data_path/init_time_reg/q_reg[0]  ( .D(n336), .CK(clk), .RN(n467), 
        .Q(curr_time[0]), .QN(n515) );
  DFFRX1 \data_path/init_time_reg/q_reg[18]  ( .D(n321), .CK(clk), .RN(n467), 
        .Q(curr_time[18]), .QN(n519) );
  DFFRX1 \data_path/init_time_reg/q_reg[23]  ( .D(n316), .CK(clk), .RN(n22), 
        .Q(curr_time[23]), .QN(n503) );
  DFFRX1 \data_path/init_time_reg/q_reg[22]  ( .D(n317), .CK(clk), .RN(n542), 
        .Q(curr_time[22]), .QN(n531) );
  DFFRX1 \data_path/init_time_reg/q_reg[21]  ( .D(n318), .CK(clk), .RN(n542), 
        .Q(curr_time[21]), .QN(n534) );
  DFFRX1 \data_path/init_time_reg/q_reg[13]  ( .D(n326), .CK(clk), .RN(n467), 
        .Q(curr_time[13]), .QN(n533) );
  DFFRX1 \data_path/init_time_reg/q_reg[3]  ( .D(n335), .CK(clk), .RN(n467), 
        .Q(curr_time[3]), .QN(n528) );
  DFFRX1 \data_path/init_time_reg/q_reg[11]  ( .D(n328), .CK(clk), .RN(n22), 
        .Q(curr_time[11]), .QN(n502) );
  DFFRX1 \data_path/so_reg/q_reg[25]  ( .D(n341), .CK(clk), .RN(n542), .Q(n777), .QN(n454) );
  DFFRX1 \data_path/so_reg/q_reg[24]  ( .D(n342), .CK(clk), .RN(n542), .Q(n778), .QN(n452) );
  DFFRX1 \data_path/so_reg/q_reg[23]  ( .D(n343), .CK(clk), .RN(n542), .Q(n779), .QN(n450) );
  DFFRX1 \data_path/so_reg/q_reg[21]  ( .D(n345), .CK(clk), .RN(n542), .Q(n781), .QN(n448) );
  DFFRX1 \data_path/so_reg/q_reg[14]  ( .D(n352), .CK(clk), .RN(n542), .Q(n783), .QN(n446) );
  DFFRX1 \data_path/so_reg/q_reg[13]  ( .D(n353), .CK(clk), .RN(n542), .Q(n784), .QN(n444) );
  DFFRX1 \data_path/so_reg/q_reg[12]  ( .D(n354), .CK(clk), .RN(n542), .Q(n785), .QN(n442) );
  DFFRX1 \data_path/so_reg/q_reg[11]  ( .D(n355), .CK(clk), .RN(n542), .Q(n786), .QN(n440) );
  DFFRX1 \data_path/so_reg/q_reg[28]  ( .D(n338), .CK(clk), .RN(n467), .Q(
        im_d_w[28]), .QN(n537) );
  DFFRX1 \data_path/so_reg/q_reg[18]  ( .D(n348), .CK(clk), .RN(n542), .Q(
        im_d_w_18), .QN(n538) );
  DFFRX1 \data_path/so_reg/q_reg[8]  ( .D(n358), .CK(clk), .RN(n542), .Q(
        im_d_w_8), .QN(n536) );
  DFFRX1 \data_path/so_reg/q_reg[26]  ( .D(n340), .CK(clk), .RN(n22), .Q(n776), 
        .QN(n456) );
  DFFRX1 \data_path/so_reg/q_reg[20]  ( .D(n346), .CK(clk), .RN(n22), .Q(n782), 
        .QN(n462) );
  DFFRX1 \data_path/so_reg/q_reg[10]  ( .D(n356), .CK(clk), .RN(n542), .Q(n787), .QN(n460) );
  DFFRX1 \data_path/so_reg/q_reg[27]  ( .D(n339), .CK(clk), .RN(n22), .Q(n775), 
        .QN(n458) );
  DFFRX1 \data_path/photo_num_reg/q_reg[0]  ( .D(n367), .CK(clk), .RN(n467), 
        .Q(photo_num[0]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[0]  ( .D(n416), .CK(clk), .RN(n22), .Q(
        fb_addr[0]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[2]  ( .D(n18), .CK(clk), .RN(n467), .Q(
        fb_addr[2]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[15]  ( .D(n383), .CK(clk), .RN(n22), .Q(
        fb_addr[15]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[14]  ( .D(n386), .CK(clk), .RN(n467), 
        .Q(fb_addr[14]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[4]  ( .D(n16), .CK(clk), .RN(n22), .Q(
        fb_addr[4]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[19]  ( .D(n374), .CK(clk), .RN(n542), 
        .Q(fb_addr[19]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[18]  ( .D(n377), .CK(clk), .RN(n542), 
        .Q(fb_addr[18]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[17]  ( .D(n380), .CK(clk), .RN(n467), 
        .Q(fb_addr[17]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[9]  ( .D(n401), .CK(clk), .RN(n542), .Q(
        fb_addr[9]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[6]  ( .D(n407), .CK(clk), .RN(n467), .Q(
        fb_addr[6]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[12]  ( .D(n392), .CK(clk), .RN(n542), 
        .Q(fb_addr[12]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[10]  ( .D(n398), .CK(clk), .RN(n22), .Q(
        fb_addr[10]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[5]  ( .D(n410), .CK(clk), .RN(n467), .Q(
        fb_addr[5]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[1]  ( .D(n20), .CK(clk), .RN(n542), .Q(
        fb_addr[1]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[8]  ( .D(n14), .CK(clk), .RN(n22), .Q(
        fb_addr[8]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[7]  ( .D(n404), .CK(clk), .RN(n542), .Q(
        fb_addr[7]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[3]  ( .D(n413), .CK(clk), .RN(n467), .Q(
        fb_addr[3]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[13]  ( .D(n389), .CK(clk), .RN(n467), 
        .Q(fb_addr[13]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[11]  ( .D(n395), .CK(clk), .RN(n22), .Q(
        fb_addr[11]) );
  DFFRX1 \data_path/fb_addr_reg/q_reg[16]  ( .D(n12), .CK(clk), .RN(n22), .Q(
        fb_addr[16]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[0]  ( .D(n415), .CK(clk), .RN(
        n22), .Q(curr_photo_addr[0]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[2]  ( .D(n17), .CK(clk), .RN(
        n467), .Q(curr_photo_addr[2]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[15]  ( .D(n382), .CK(clk), .RN(
        n22), .Q(curr_photo_addr[15]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[14]  ( .D(n385), .CK(clk), .RN(
        n467), .Q(curr_photo_addr[14]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[4]  ( .D(n15), .CK(clk), .RN(n22), .Q(curr_photo_addr[4]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[19]  ( .D(n373), .CK(clk), .RN(
        n542), .Q(curr_photo_addr[19]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[18]  ( .D(n376), .CK(clk), .RN(
        n467), .Q(curr_photo_addr[18]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[17]  ( .D(n379), .CK(clk), .RN(
        n467), .Q(curr_photo_addr[17]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[9]  ( .D(n400), .CK(clk), .RN(
        n542), .Q(curr_photo_addr[9]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[6]  ( .D(n406), .CK(clk), .RN(
        n467), .Q(curr_photo_addr[6]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[12]  ( .D(n391), .CK(clk), .RN(
        n467), .Q(curr_photo_addr[12]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[10]  ( .D(n397), .CK(clk), .RN(
        n542), .Q(curr_photo_addr[10]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[5]  ( .D(n409), .CK(clk), .RN(
        n467), .Q(curr_photo_addr[5]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[1]  ( .D(n19), .CK(clk), .RN(
        n467), .Q(curr_photo_addr[1]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[8]  ( .D(n13), .CK(clk), .RN(n22), .Q(curr_photo_addr[8]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[7]  ( .D(n403), .CK(clk), .RN(
        n542), .Q(curr_photo_addr[7]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[3]  ( .D(n412), .CK(clk), .RN(
        n467), .Q(curr_photo_addr[3]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[13]  ( .D(n388), .CK(clk), .RN(
        n467), .Q(curr_photo_addr[13]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[11]  ( .D(n394), .CK(clk), .RN(
        n22), .Q(curr_photo_addr[11]) );
  DFFRX1 \data_path/curr_photo_addr_reg/q_reg[16]  ( .D(n11), .CK(clk), .RN(
        n22), .Q(curr_photo_addr[16]) );
  DFFRX1 \data_path/init_time_reg/q_reg[20]  ( .D(n319), .CK(clk), .RN(n542), 
        .Q(curr_time[20]) );
  DFFRX1 \data_path/init_time_reg/q_reg[5]  ( .D(n334), .CK(clk), .RN(n467), 
        .Q(curr_time[5]) );
  DFFRX1 \data_path/init_time_reg/q_reg[8]  ( .D(n331), .CK(clk), .RN(n22), 
        .Q(curr_time[8]) );
  DFFRX1 \data_path/so_reg/q_reg[29]  ( .D(n337), .CK(clk), .RN(n542), .Q(
        im_d_w[29]) );
  DFFRX1 \data_path/so_reg/q_reg[19]  ( .D(n347), .CK(clk), .RN(n467), .Q(
        im_d_w_19) );
  DFFRX1 \data_path/so_reg/q_reg[9]  ( .D(n357), .CK(clk), .RN(n467), .Q(
        im_d_w_9) );
  DFFRX1 \data_path/so_reg/q_reg[1]  ( .D(n365), .CK(clk), .RN(n467), .QN(n477) );
  DFFRX1 \data_path/so_reg/q_reg[15]  ( .D(n351), .CK(clk), .RN(n467), .QN(
        n484) );
  DFFRX1 \data_path/so_reg/q_reg[5]  ( .D(n361), .CK(clk), .RN(n467), .QN(n488) );
  DFFRX1 \data_path/so_reg/q_reg[22]  ( .D(n344), .CK(clk), .RN(n467), .Q(n780) );
  DFFRX1 \data_path/so_reg/q_reg[4]  ( .D(n362), .CK(clk), .RN(n467), .QN(n486) );
  DFFRX1 \data_path/so_reg/q_reg[3]  ( .D(n363), .CK(clk), .RN(n467), .QN(n482) );
  DFFRX1 \data_path/so_reg/q_reg[2]  ( .D(n364), .CK(clk), .RN(n467), .QN(n480) );
  DFFRX1 \data_path/so_reg/q_reg[16]  ( .D(n350), .CK(clk), .RN(n467), .QN(
        n473) );
  DFFRX1 \data_path/so_reg/q_reg[6]  ( .D(n360), .CK(clk), .RN(n467), .QN(n490) );
  DFFRX1 \data_path/so_reg/q_reg[0]  ( .D(n366), .CK(clk), .RN(n467), .QN(n475) );
  DFFRX1 \data_path/so_reg/q_reg[17]  ( .D(n349), .CK(clk), .RN(n467), .QN(
        n492) );
  DFFRX1 \data_path/so_reg/q_reg[7]  ( .D(n359), .CK(clk), .RN(n467), .QN(n494) );
  AND2X2 U435 ( .A(si_sel), .B(en_si), .Y(n717) );
  INVX4 U436 ( .A(en_si), .Y(n731) );
  BUFX8 U437 ( .A(n542), .Y(n467) );
  INVX8 U438 ( .A(reset), .Y(n22) );
  CLKBUFX8 U439 ( .A(n22), .Y(n542) );
  NOR4X1 U440 ( .A(\data_path/si_w[16] ), .B(\data_path/si_w[17] ), .C(
        \data_path/si_w[18] ), .D(\data_path/si_w[19] ), .Y(n421) );
  NOR4X1 U441 ( .A(\data_path/si_w[1] ), .B(\data_path/si_w[2] ), .C(
        \data_path/si_w[15] ), .D(\data_path/si_w[23] ), .Y(n422) );
  NOR4X1 U442 ( .A(\data_path/si_w[20] ), .B(\data_path/si_w[14] ), .C(
        \data_path/si_w[21] ), .D(\data_path/si_w[22] ), .Y(n423) );
  AND4X1 U443 ( .A(n422), .B(n423), .C(n520), .D(en_curr_photo_size), .Y(n424)
         );
  AND4X1 U444 ( .A(n500), .B(n421), .C(n507), .D(n424), .Y(n548) );
  AO22X1 U445 ( .A0(n539), .A1(\intadd_1/SUM[2] ), .B0(\intadd_1/SUM[1] ), 
        .B1(n540), .Y(n425) );
  AOI211X1 U446 ( .A0(n727), .A1(n786), .B0(n634), .C0(n425), .Y(n426) );
  NAND2X1 U447 ( .A(\intadd_1/SUM[0] ), .B(n640), .Y(n427) );
  OAI211X1 U448 ( .A0(n466), .A1(n521), .B0(n426), .C0(n427), .Y(n355) );
  AO22X1 U449 ( .A0(n539), .A1(\intadd_1/SUM[3] ), .B0(\intadd_1/SUM[2] ), 
        .B1(n540), .Y(n428) );
  AOI211X1 U450 ( .A0(n727), .A1(n785), .B0(n634), .C0(n428), .Y(n429) );
  NAND2XL U451 ( .A(\intadd_1/SUM[1] ), .B(n640), .Y(n430) );
  OAI211X1 U452 ( .A0(n466), .A1(n499), .B0(n429), .C0(n430), .Y(n354) );
  AO22X1 U453 ( .A0(n539), .A1(\intadd_1/SUM[4] ), .B0(\intadd_1/SUM[3] ), 
        .B1(n540), .Y(n431) );
  AOI211X1 U454 ( .A0(n727), .A1(n784), .B0(n634), .C0(n431), .Y(n432) );
  NAND2XL U455 ( .A(\intadd_1/SUM[2] ), .B(n640), .Y(n433) );
  OAI211X1 U456 ( .A0(n466), .A1(n501), .B0(n432), .C0(n433), .Y(n353) );
  AO22X1 U457 ( .A0(n539), .A1(\intadd_1/SUM[5] ), .B0(\intadd_1/SUM[4] ), 
        .B1(n540), .Y(n434) );
  AOI211X1 U458 ( .A0(n727), .A1(n783), .B0(n634), .C0(n434), .Y(n435) );
  NAND2XL U459 ( .A(\intadd_1/SUM[3] ), .B(n640), .Y(n436) );
  OAI211X1 U460 ( .A0(n466), .A1(n520), .B0(n435), .C0(n436), .Y(n352) );
  AO22X1 U461 ( .A0(n539), .A1(\intadd_0/SUM[2] ), .B0(\intadd_0/SUM[1] ), 
        .B1(n540), .Y(n437) );
  AOI211X1 U462 ( .A0(n727), .A1(n781), .B0(n634), .C0(n437), .Y(n438) );
  NAND2X1 U463 ( .A(\intadd_0/SUM[0] ), .B(n640), .Y(n439) );
  OAI211X1 U464 ( .A0(n466), .A1(n525), .B0(n438), .C0(n439), .Y(n345) );
  AOI211X1 U465 ( .A0(curr_time[13]), .A1(n669), .B0(curr_time[15]), .C0(
        curr_time[14]), .Y(n676) );
  INVX16 U466 ( .A(n440), .Y(IM_D[9]) );
  INVX16 U467 ( .A(n442), .Y(IM_D[10]) );
  INVX16 U468 ( .A(n444), .Y(IM_D[11]) );
  INVX16 U469 ( .A(n446), .Y(IM_D[12]) );
  INVX16 U470 ( .A(n448), .Y(IM_D[17]) );
  INVX16 U471 ( .A(n450), .Y(IM_D[19]) );
  INVX16 U472 ( .A(n452), .Y(IM_D[20]) );
  INVX16 U473 ( .A(n454), .Y(IM_D[21]) );
  INVX16 U474 ( .A(n456), .Y(IM_D[22]) );
  INVX16 U475 ( .A(n458), .Y(IM_D[23]) );
  INVX16 U476 ( .A(n460), .Y(IM_D[8]) );
  INVX16 U477 ( .A(n462), .Y(IM_D[16]) );
  INVX8 U478 ( .A(n544), .Y(n464) );
  INVX8 U479 ( .A(n543), .Y(n465) );
  BUFX4 U480 ( .A(n641), .Y(n466) );
  NOR2X1 U481 ( .A(n657), .B(n659), .Y(n665) );
  AOI211X1 U482 ( .A0(n470), .A1(n654), .B0(n670), .C0(n663), .Y(n655) );
  BUFX4 U483 ( .A(n730), .Y(n541) );
  INVX6 U484 ( .A(en_so), .Y(n727) );
  OA21XL U485 ( .A0(IM_D[0]), .A1(n728), .B0(n466), .Y(n555) );
  OA21XL U486 ( .A0(\data_path/si_w[0] ), .A1(n615), .B0(en_so), .Y(n554) );
  NOR2X6 U487 ( .A(n727), .B(n615), .Y(n640) );
  INVX1 U488 ( .A(n468), .Y(n544) );
  INVX1 U489 ( .A(n469), .Y(n543) );
  AOI211X1 U490 ( .A0(n688), .A1(curr_time[20]), .B0(n676), .C0(n675), .Y(n678) );
  INVX16 U491 ( .A(n484), .Y(IM_D[13]) );
  BUFX16 U492 ( .A(n780), .Y(IM_D[18]) );
  NAND2X1 U493 ( .A(n710), .B(n709), .Y(n719) );
  NOR2X1 U494 ( .A(n505), .B(n708), .Y(n709) );
  NOR2X1 U495 ( .A(n528), .B(n657), .Y(n660) );
  NAND2X1 U496 ( .A(n470), .B(n654), .Y(n657) );
  NOR2X1 U497 ( .A(n699), .B(n723), .Y(n703) );
  NOR2X1 U498 ( .A(curr_time[8]), .B(n714), .Y(n699) );
  CLKINVX1 U499 ( .A(n648), .Y(n659) );
  NOR2X1 U500 ( .A(n670), .B(n663), .Y(n648) );
  NOR2X1 U501 ( .A(n506), .B(n686), .Y(n681) );
  NAND2X1 U502 ( .A(en_init_time), .B(n678), .Y(n686) );
  AOI211X1 U503 ( .A0(n646), .A1(curr_time[5]), .B0(curr_time[6]), .C0(
        curr_time[7]), .Y(n668) );
  OAI21X1 U504 ( .A0(curr_time[16]), .A1(n687), .B0(n721), .Y(n682) );
  CLKINVX1 U505 ( .A(n678), .Y(n687) );
  OAI21X1 U506 ( .A0(n688), .A1(n687), .B0(n721), .Y(n691) );
  NOR2BX1 U507 ( .AN(n688), .B(n686), .Y(n690) );
  NOR3X2 U508 ( .A(n679), .B(n506), .C(n519), .Y(n688) );
  OAI21X1 U509 ( .A0(\intadd_0/n1 ), .A1(im_d_w[28]), .B0(n638), .Y(n693) );
  NAND2X1 U510 ( .A(\intadd_0/n1 ), .B(im_d_w[28]), .Y(n638) );
  OAI31X1 U511 ( .A0(n560), .A1(n559), .A2(n558), .B0(expand_sel[3]), .Y(n574)
         );
  NOR2X1 U512 ( .A(n470), .B(n654), .Y(n652) );
  NOR2X2 U513 ( .A(n649), .B(n515), .Y(n654) );
  CLKINVX1 U514 ( .A(n539), .Y(n639) );
  BUFX4 U515 ( .A(n629), .Y(n539) );
  BUFX4 U516 ( .A(n635), .Y(n540) );
  NOR2X1 U517 ( .A(si_sel), .B(n731), .Y(n730) );
  INVX16 U518 ( .A(n774), .Y(IM_A[0]) );
  INVX16 U519 ( .A(n773), .Y(IM_A[1]) );
  INVX16 U520 ( .A(n772), .Y(IM_A[2]) );
  INVX16 U521 ( .A(n771), .Y(IM_A[3]) );
  INVX16 U522 ( .A(n770), .Y(IM_A[4]) );
  INVX16 U523 ( .A(n769), .Y(IM_A[5]) );
  INVX16 U524 ( .A(n768), .Y(IM_A[6]) );
  INVX16 U525 ( .A(n767), .Y(IM_A[7]) );
  INVX16 U526 ( .A(n766), .Y(IM_A[8]) );
  INVX16 U527 ( .A(n765), .Y(IM_A[9]) );
  INVX16 U528 ( .A(n764), .Y(IM_A[10]) );
  INVX16 U529 ( .A(n763), .Y(IM_A[11]) );
  INVX16 U530 ( .A(n762), .Y(IM_A[12]) );
  INVX16 U531 ( .A(n761), .Y(IM_A[13]) );
  INVX16 U532 ( .A(n760), .Y(IM_A[14]) );
  INVX16 U533 ( .A(n759), .Y(IM_A[15]) );
  INVX16 U534 ( .A(n758), .Y(IM_A[16]) );
  INVX16 U535 ( .A(n757), .Y(IM_A[17]) );
  INVX16 U536 ( .A(n756), .Y(IM_A[18]) );
  CLKINVX1 U537 ( .A(n754), .Y(n471) );
  INVX16 U538 ( .A(n471), .Y(IM_A[19]) );
  INVX16 U539 ( .A(n473), .Y(IM_D[14]) );
  INVX16 U540 ( .A(n475), .Y(IM_D[0]) );
  INVX16 U541 ( .A(n477), .Y(IM_D[1]) );
  INVX16 U542 ( .A(n480), .Y(IM_D[2]) );
  INVX16 U543 ( .A(n482), .Y(IM_D[3]) );
  INVX16 U544 ( .A(n486), .Y(IM_D[4]) );
  INVX16 U545 ( .A(n488), .Y(IM_D[5]) );
  INVX16 U546 ( .A(n490), .Y(IM_D[6]) );
  INVX16 U547 ( .A(n492), .Y(IM_D[15]) );
  INVX16 U548 ( .A(n494), .Y(IM_D[7]) );
  OAI21X1 U549 ( .A0(\intadd_2/n1 ), .A1(im_d_w_8), .B0(n596), .Y(n600) );
  NAND2X1 U550 ( .A(\intadd_2/n1 ), .B(im_d_w_8), .Y(n596) );
  OAI21X1 U551 ( .A0(\intadd_1/n1 ), .A1(im_d_w_18), .B0(n611), .Y(n725) );
  NAND2X1 U552 ( .A(\intadd_1/n1 ), .B(im_d_w_18), .Y(n611) );
  NOR2X1 U553 ( .A(\data_path/si_w[4] ), .B(n546), .Y(n549) );
  NAND4X1 U554 ( .A(n499), .B(n501), .C(n508), .D(n522), .Y(n546) );
  NOR2BX1 U555 ( .AN(init_time_mux_sel), .B(n668), .Y(n674) );
  NAND2X1 U556 ( .A(n668), .B(init_time_mux_sel), .Y(n663) );
  CLKINVX1 U557 ( .A(n710), .Y(n714) );
  NOR2X1 U558 ( .A(n672), .B(n670), .Y(n710) );
  NAND2X1 U559 ( .A(expand_sel[0]), .B(n566), .Y(n567) );
  CLKINVX1 U560 ( .A(expand_sel[1]), .Y(n566) );
  NAND2X1 U561 ( .A(n553), .B(so_mux_sel[0]), .Y(n615) );
  NAND2XL U562 ( .A(IM_D[14]), .B(n727), .Y(n609) );
  NOR2X1 U563 ( .A(n496), .B(n497), .Y(n576) );
  NOR2X1 U564 ( .A(n555), .B(n498), .Y(n496) );
  NOR2XL U565 ( .A(n554), .B(n475), .Y(n497) );
  NOR2X2 U566 ( .A(expand_sel[1]), .B(expand_sel[0]), .Y(n569) );
  INVX3 U567 ( .A(n640), .Y(n728) );
  INVX3 U568 ( .A(n724), .Y(n722) );
  NOR2X4 U569 ( .A(init_time_mux_sel), .B(n670), .Y(n724) );
  INVX4 U570 ( .A(n644), .Y(n634) );
  NAND4X2 U571 ( .A(so_mux_sel[1]), .B(n575), .C(n574), .D(n573), .Y(n644) );
  NOR2BX2 U572 ( .AN(n672), .B(n723), .Y(n721) );
  NAND2X2 U573 ( .A(en_init_time), .B(n663), .Y(n723) );
  NAND2XL U574 ( .A(n776), .B(n727), .Y(n636) );
  AOI211XL U575 ( .A0(n775), .A1(n727), .B0(n643), .C0(n642), .Y(n645) );
  AOI22XL U576 ( .A0(\data_path/si_w[8] ), .A1(n602), .B0(n787), .B1(n601), 
        .Y(n603) );
  AOI22XL U577 ( .A0(\data_path/si_w[16] ), .A1(n617), .B0(n782), .B1(n616), 
        .Y(n618) );
  INVXL U578 ( .A(n707), .Y(n399) );
  INVXL U579 ( .A(n545), .Y(n417) );
  INVXL U580 ( .A(n712), .Y(n396) );
  INVXL U581 ( .A(n696), .Y(n411) );
  INVXL U582 ( .A(n695), .Y(n414) );
  INVXL U583 ( .A(n698), .Y(n405) );
  INVXL U584 ( .A(n697), .Y(n408) );
  INVXL U585 ( .A(n718), .Y(n393) );
  INVXL U586 ( .A(n702), .Y(n402) );
  INVXL U587 ( .A(en_photo_num), .Y(n733) );
  OAI211XL U588 ( .A0(en_curr_photo_size), .A1(n514), .B0(n551), .C0(n734), 
        .Y(n368) );
  NAND4XL U589 ( .A(\data_path/si_w[7] ), .B(n549), .C(n548), .D(n547), .Y(
        n551) );
  NOR3XL U590 ( .A(\data_path/si_w[9] ), .B(\data_path/si_w[0] ), .C(
        \data_path/si_w[3] ), .Y(n547) );
  NAND4XL U591 ( .A(n550), .B(n549), .C(n548), .D(n517), .Y(n734) );
  INVXL U592 ( .A(n652), .Y(n653) );
  AOI211XL U593 ( .A0(curr_time[4]), .A1(n670), .B0(n662), .C0(n661), .Y(n141)
         );
  NOR2XL U594 ( .A(n722), .B(n509), .Y(n661) );
  AOI211XL U595 ( .A0(curr_time[4]), .A1(n660), .B0(n659), .C0(n658), .Y(n662)
         );
  NOR2XL U596 ( .A(curr_time[4]), .B(n660), .Y(n658) );
  NOR2XL U597 ( .A(n651), .B(n650), .Y(n145) );
  AOI211XL U598 ( .A0(n649), .A1(n515), .B0(n654), .C0(n659), .Y(n651) );
  INVXL U599 ( .A(n667), .Y(n334) );
  INVXL U600 ( .A(n664), .Y(n666) );
  OAI32XL U601 ( .A0(n528), .A1(n655), .A2(n670), .B0(n665), .B1(curr_time[3]), 
        .Y(n656) );
  NAND2XL U602 ( .A(curr_time[12]), .B(curr_time[11]), .Y(n720) );
  AOI21XL U603 ( .A0(curr_time[8]), .A1(n723), .B0(n699), .Y(n671) );
  AOI22XL U604 ( .A0(curr_time[12]), .A1(n715), .B0(n724), .B1(
        \data_path/si_w[12] ), .Y(n716) );
  AOI22XL U605 ( .A0(curr_time[10]), .A1(n704), .B0(\data_path/si_w[10] ), 
        .B1(n724), .Y(n705) );
  NAND2XL U606 ( .A(curr_time[8]), .B(n710), .Y(n706) );
  OAI211XL U607 ( .A0(n722), .A1(n524), .B0(n685), .C0(n684), .Y(n321) );
  NOR2XL U608 ( .A(n687), .B(curr_time[17]), .Y(n683) );
  NAND3XL U609 ( .A(curr_time[17]), .B(n681), .C(n519), .Y(n685) );
  INVXL U610 ( .A(n692), .Y(n319) );
  NAND2XL U611 ( .A(n674), .B(n676), .Y(n672) );
  NAND3XL U612 ( .A(n674), .B(n673), .C(n503), .Y(n675) );
  AOI211XL U613 ( .A0(curr_time[20]), .A1(curr_time[19]), .B0(curr_time[21]), 
        .C0(curr_time[22]), .Y(n673) );
  NOR2XL U614 ( .A(n652), .B(n664), .Y(n646) );
  NAND2XL U615 ( .A(curr_time[4]), .B(curr_time[3]), .Y(n664) );
  AOI211XL U616 ( .A0(n505), .A1(n708), .B0(n518), .C0(n502), .Y(n669) );
  NAND2XL U617 ( .A(curr_time[9]), .B(curr_time[8]), .Y(n708) );
  CLKINVX2 U618 ( .A(en_init_time), .Y(n670) );
  OAI211XL U619 ( .A0(n466), .A1(n516), .B0(n586), .C0(n585), .Y(n363) );
  NAND2XL U620 ( .A(n640), .B(\intadd_2/SUM[2] ), .Y(n585) );
  AOI211XL U621 ( .A0(n540), .A1(\intadd_2/SUM[3] ), .B0(n634), .C0(n584), .Y(
        n586) );
  OAI211XL U622 ( .A0(n466), .A1(n509), .B0(n589), .C0(n588), .Y(n362) );
  NAND2XL U623 ( .A(n640), .B(\intadd_2/SUM[3] ), .Y(n588) );
  AOI211XL U624 ( .A0(n540), .A1(\intadd_2/SUM[4] ), .B0(n634), .C0(n587), .Y(
        n589) );
  OAI211XL U625 ( .A0(n466), .A1(n526), .B0(n625), .C0(n624), .Y(n343) );
  NAND2XL U626 ( .A(n640), .B(\intadd_0/SUM[2] ), .Y(n624) );
  AOI211XL U627 ( .A0(n540), .A1(\intadd_0/SUM[3] ), .B0(n634), .C0(n623), .Y(
        n625) );
  OAI211XL U628 ( .A0(n466), .A1(n504), .B0(n580), .C0(n579), .Y(n365) );
  NAND2XL U629 ( .A(n640), .B(\intadd_2/SUM[0] ), .Y(n579) );
  AOI211XL U630 ( .A0(\intadd_2/SUM[1] ), .A1(n540), .B0(n634), .C0(n578), .Y(
        n580) );
  OAI211XL U631 ( .A0(n466), .A1(n532), .B0(n628), .C0(n627), .Y(n342) );
  NAND2XL U632 ( .A(n640), .B(\intadd_0/SUM[3] ), .Y(n627) );
  AOI211XL U633 ( .A0(n540), .A1(\intadd_0/SUM[4] ), .B0(n634), .C0(n626), .Y(
        n628) );
  OAI211XL U634 ( .A0(n466), .A1(n510), .B0(n583), .C0(n582), .Y(n364) );
  NAND2XL U635 ( .A(n640), .B(\intadd_2/SUM[1] ), .Y(n582) );
  AOI211XL U636 ( .A0(n540), .A1(\intadd_2/SUM[2] ), .B0(n634), .C0(n581), .Y(
        n583) );
  OAI211XL U637 ( .A0(n507), .A1(n466), .B0(n607), .C0(n606), .Y(n351) );
  NAND2XL U638 ( .A(n640), .B(\intadd_1/SUM[4] ), .Y(n606) );
  AOI211XL U639 ( .A0(n540), .A1(\intadd_1/SUM[5] ), .B0(n634), .C0(n605), .Y(
        n607) );
  OAI211XL U640 ( .A0(n466), .A1(n524), .B0(n622), .C0(n621), .Y(n344) );
  NAND2XL U641 ( .A(n640), .B(\intadd_0/SUM[1] ), .Y(n621) );
  AOI211XL U642 ( .A0(n540), .A1(\intadd_0/SUM[2] ), .B0(n634), .C0(n620), .Y(
        n622) );
  OAI211XL U643 ( .A0(n466), .A1(n508), .B0(n592), .C0(n591), .Y(n361) );
  NAND2XL U644 ( .A(n640), .B(\intadd_2/SUM[4] ), .Y(n591) );
  AOI211XL U645 ( .A0(n540), .A1(\intadd_2/SUM[5] ), .B0(n634), .C0(n590), .Y(
        n592) );
  OAI211XL U646 ( .A0(n511), .A1(n466), .B0(n632), .C0(n631), .Y(n341) );
  NAND2XL U647 ( .A(n640), .B(\intadd_0/SUM[4] ), .Y(n631) );
  AOI211XL U648 ( .A0(n540), .A1(\intadd_0/SUM[5] ), .B0(n634), .C0(n630), .Y(
        n632) );
  OAI211XL U649 ( .A0(n693), .A1(n639), .B0(n637), .C0(n636), .Y(n340) );
  AOI211XL U650 ( .A0(n540), .A1(\intadd_0/SUM[6] ), .B0(n634), .C0(n633), .Y(
        n637) );
  OAI211XL U651 ( .A0(n600), .A1(n639), .B0(n595), .C0(n594), .Y(n360) );
  NAND2X1 U652 ( .A(IM_D[6]), .B(n727), .Y(n594) );
  AOI211XL U653 ( .A0(n540), .A1(\intadd_2/SUM[6] ), .B0(n634), .C0(n593), .Y(
        n595) );
  OAI211XL U654 ( .A0(n725), .A1(n639), .B0(n610), .C0(n609), .Y(n350) );
  AOI211XL U655 ( .A0(n540), .A1(\intadd_1/SUM[6] ), .B0(n634), .C0(n608), .Y(
        n610) );
  OAI211XL U656 ( .A0(n726), .A1(n693), .B0(n645), .C0(n644), .Y(n339) );
  NOR2XL U657 ( .A(n639), .B(n694), .Y(n643) );
  OAI211XL U658 ( .A0(n726), .A1(n725), .B0(n614), .C0(n644), .Y(n349) );
  AOI211X1 U659 ( .A0(IM_D[15]), .A1(n727), .B0(n613), .C0(n612), .Y(n614) );
  NOR2XL U660 ( .A(n639), .B(n729), .Y(n613) );
  OAI211XL U661 ( .A0(n726), .A1(n600), .B0(n599), .C0(n644), .Y(n359) );
  AOI211X1 U662 ( .A0(IM_D[7]), .A1(n727), .B0(n598), .C0(n597), .Y(n599) );
  NOR2XL U663 ( .A(n639), .B(n701), .Y(n598) );
  NAND3XL U664 ( .A(n577), .B(n576), .C(n644), .Y(n366) );
  AOI22XL U665 ( .A0(n539), .A1(\intadd_2/SUM[1] ), .B0(n540), .B1(
        \intadd_2/SUM[0] ), .Y(n577) );
  NOR2BXL U666 ( .AN(IM_D[0]), .B(n498), .Y(\intadd_2/CI ) );
  NAND3XL U667 ( .A(n619), .B(n618), .C(n644), .Y(n346) );
  OAI21XL U668 ( .A0(n782), .A1(n728), .B0(n466), .Y(n617) );
  AOI22XL U669 ( .A0(n539), .A1(\intadd_0/SUM[1] ), .B0(n540), .B1(
        \intadd_0/SUM[0] ), .Y(n619) );
  AND2XL U670 ( .A(\data_path/si_w[16] ), .B(n782), .Y(\intadd_0/CI ) );
  NAND3XL U671 ( .A(n604), .B(n603), .C(n644), .Y(n356) );
  INVXL U672 ( .A(expand_sel[3]), .Y(n570) );
  AOI211XL U673 ( .A0(n569), .A1(\data_path/si_w[12] ), .B0(expand_sel[2]), 
        .C0(n568), .Y(n571) );
  AOI211XL U674 ( .A0(n569), .A1(\data_path/si_w[8] ), .B0(n563), .C0(n562), 
        .Y(n572) );
  AOI211XL U675 ( .A0(n569), .A1(\data_path/si_w[4] ), .B0(expand_sel[2]), 
        .C0(n557), .Y(n558) );
  INVXL U676 ( .A(expand_sel[0]), .Y(n564) );
  NOR2XL U677 ( .A(\data_path/si_w[0] ), .B(n563), .Y(n559) );
  NOR2XL U678 ( .A(n569), .B(n563), .Y(n560) );
  INVXL U679 ( .A(expand_sel[2]), .Y(n563) );
  NOR2XL U680 ( .A(so_mux_sel[0]), .B(n727), .Y(n575) );
  OAI21XL U681 ( .A0(n787), .A1(n728), .B0(n466), .Y(n602) );
  INVXL U682 ( .A(so_mux_sel[1]), .Y(n553) );
  AOI22XL U683 ( .A0(n539), .A1(\intadd_1/SUM[1] ), .B0(n540), .B1(
        \intadd_1/SUM[0] ), .Y(n604) );
  NOR2BXL U684 ( .AN(n787), .B(n500), .Y(\intadd_1/CI ) );
  NOR2BXL U685 ( .AN(\sftr_n[0] ), .B(n552), .Y(n629) );
  NAND3XL U686 ( .A(so_mux_sel[1]), .B(so_mux_sel[0]), .C(en_so), .Y(n552) );
  INVXL U687 ( .A(n755), .Y(n754) );
  AOI222XL U688 ( .A0(n731), .A1(\data_path/si_w[2] ), .B0(n541), .B1(IM_Q[2]), 
        .C0(n717), .C1(CR_Q[2]), .Y(n314) );
  AOI222XL U689 ( .A0(n731), .A1(\data_path/si_w[4] ), .B0(n541), .B1(IM_Q[4]), 
        .C0(n717), .C1(CR_Q[4]), .Y(n313) );
  AOI222XL U690 ( .A0(n731), .A1(\data_path/si_w[8] ), .B0(n541), .B1(IM_Q[8]), 
        .C0(n717), .C1(CR_Q[8]), .Y(n312) );
  AOI222XL U691 ( .A0(n731), .A1(\data_path/si_w[1] ), .B0(n717), .B1(CR_Q[1]), 
        .C0(IM_Q[1]), .C1(n541), .Y(n315) );
  AOI222XL U692 ( .A0(n731), .A1(\data_path/si_w[10] ), .B0(n541), .B1(
        IM_Q[10]), .C0(n717), .C1(CR_Q[10]), .Y(n707) );
  AOI222XL U693 ( .A0(n731), .A1(\data_path/si_w[0] ), .B0(n541), .B1(IM_Q[0]), 
        .C0(n717), .C1(CR_Q[0]), .Y(n545) );
  AOI222XL U694 ( .A0(n731), .A1(\data_path/si_w[11] ), .B0(n541), .B1(
        IM_Q[11]), .C0(n717), .C1(CR_Q[11]), .Y(n712) );
  AOI222XL U695 ( .A0(n731), .A1(\data_path/si_w[5] ), .B0(n541), .B1(IM_Q[5]), 
        .C0(n717), .C1(CR_Q[5]), .Y(n696) );
  AOI222XL U696 ( .A0(n731), .A1(\data_path/si_w[3] ), .B0(n541), .B1(IM_Q[3]), 
        .C0(n717), .C1(CR_Q[3]), .Y(n695) );
  AOI222XL U697 ( .A0(n731), .A1(\data_path/si_w[7] ), .B0(n541), .B1(IM_Q[7]), 
        .C0(n717), .C1(CR_Q[7]), .Y(n698) );
  AOI222XL U698 ( .A0(n731), .A1(\data_path/si_w[6] ), .B0(n541), .B1(IM_Q[6]), 
        .C0(n717), .C1(CR_Q[6]), .Y(n697) );
  AOI222XL U699 ( .A0(n731), .A1(\data_path/si_w[12] ), .B0(n541), .B1(
        IM_Q[12]), .C0(n717), .C1(CR_Q[12]), .Y(n718) );
  AOI222XL U700 ( .A0(n731), .A1(\data_path/si_w[9] ), .B0(n541), .B1(IM_Q[9]), 
        .C0(n717), .C1(CR_Q[9]), .Y(n702) );
  OAI22XL U701 ( .A0(en_photo_num), .A1(n10), .B0(n733), .B1(n732), .Y(n21) );
  NOR3XL U702 ( .A(\data_path/si_w[0] ), .B(\data_path/si_w[3] ), .C(n521), 
        .Y(n550) );
  AOI222XL U703 ( .A0(n670), .A1(n470), .B0(n724), .B1(\data_path/si_w[2] ), 
        .C0(n653), .C1(n655), .Y(n144) );
  AOI222XL U704 ( .A0(\data_path/si_w[5] ), .A1(n724), .B0(curr_time[5]), .B1(
        n723), .C0(n666), .C1(n665), .Y(n667) );
  OAI222XL U705 ( .A0(n507), .A1(n722), .B0(n533), .B1(n721), .C0(n720), .C1(
        n719), .Y(n326) );
  OAI21XL U706 ( .A0(n713), .A1(n502), .B0(n711), .Y(n328) );
  OAI31XL U707 ( .A0(curr_time[12]), .A1(n502), .A2(n719), .B0(n716), .Y(n327)
         );
  OAI31XL U708 ( .A0(curr_time[10]), .A1(n529), .A2(n706), .B0(n705), .Y(n329)
         );
  AOI222XL U709 ( .A0(n691), .A1(curr_time[20]), .B0(curr_time[19]), .B1(n690), 
        .C0(n724), .C1(\data_path/si_w[20] ), .Y(n692) );
  OAI2BB2XL U710 ( .B0(n729), .B1(n728), .A0N(im_d_w_19), .A1N(n727), .Y(n347)
         );
  OAI2BB2XL U711 ( .B0(n694), .B1(n728), .A0N(im_d_w[29]), .A1N(n727), .Y(n337) );
  OAI2BB2XL U712 ( .B0(n701), .B1(n728), .A0N(im_d_w_9), .A1N(n727), .Y(n357)
         );
  OAI222XL U713 ( .A0(n701), .A1(n726), .B0(n536), .B1(en_so), .C0(n600), .C1(
        n728), .Y(n358) );
  OAI222XL U714 ( .A0(n694), .A1(n726), .B0(n537), .B1(en_so), .C0(n693), .C1(
        n728), .Y(n338) );
  OAI222XL U715 ( .A0(n729), .A1(n726), .B0(n538), .B1(en_so), .C0(n725), .C1(
        n728), .Y(n348) );
  CLKINVX1 U716 ( .A(n540), .Y(n726) );
  NOR2X1 U717 ( .A(\sftr_n[0] ), .B(n552), .Y(n635) );
  AO22X1 U718 ( .A0(\data_path/si_w[16] ), .A1(n731), .B0(n541), .B1(IM_Q[16]), 
        .Y(n418) );
  AOI2BB2X1 U719 ( .B0(n464), .B1(n498), .A0N(n464), .A1N(fb_addr[0]), .Y(n416) );
  AOI2BB2X1 U720 ( .B0(n465), .B1(n498), .A0N(n465), .A1N(curr_photo_addr[0]), 
        .Y(n415) );
  AOI2BB2X1 U721 ( .B0(n464), .B1(n516), .A0N(n464), .A1N(fb_addr[3]), .Y(n413) );
  AOI2BB2X1 U722 ( .B0(n465), .B1(n516), .A0N(n465), .A1N(curr_photo_addr[3]), 
        .Y(n412) );
  AOI2BB2X1 U723 ( .B0(n464), .B1(n508), .A0N(n464), .A1N(fb_addr[5]), .Y(n410) );
  AOI2BB2X1 U724 ( .B0(n465), .B1(n508), .A0N(n465), .A1N(curr_photo_addr[5]), 
        .Y(n409) );
  AOI2BB2X1 U725 ( .B0(n464), .B1(n522), .A0N(n464), .A1N(fb_addr[6]), .Y(n407) );
  AOI2BB2X1 U726 ( .B0(n465), .B1(n522), .A0N(n465), .A1N(curr_photo_addr[6]), 
        .Y(n406) );
  AOI2BB2X1 U727 ( .B0(n464), .B1(n517), .A0N(n464), .A1N(fb_addr[7]), .Y(n404) );
  AOI2BB2X1 U728 ( .B0(n465), .B1(n517), .A0N(n465), .A1N(curr_photo_addr[7]), 
        .Y(n403) );
  AOI2BB2X1 U729 ( .B0(en_photo_num), .B1(\data_path/si_w[0] ), .A0N(
        en_photo_num), .A1N(photo_num[0]), .Y(n367) );
  NAND3BX1 U730 ( .AN(so_mux_sel[0]), .B(en_so), .C(n553), .Y(n641) );
  OAI22XL U731 ( .A0(expand_sel[0]), .A1(\data_path/si_w[2] ), .B0(n564), .B1(
        \data_path/si_w[1] ), .Y(n556) );
  OAI22XL U732 ( .A0(n566), .A1(n556), .B0(n516), .B1(n567), .Y(n557) );
  OAI22XL U733 ( .A0(expand_sel[0]), .A1(\data_path/si_w[6] ), .B0(n564), .B1(
        \data_path/si_w[5] ), .Y(n561) );
  OAI22XL U734 ( .A0(n566), .A1(n561), .B0(n567), .B1(n517), .Y(n562) );
  OAI22XL U735 ( .A0(expand_sel[0]), .A1(\data_path/si_w[10] ), .B0(n564), 
        .B1(\data_path/si_w[9] ), .Y(n565) );
  OAI22XL U736 ( .A0(n501), .A1(n567), .B0(n566), .B1(n565), .Y(n568) );
  OAI21XL U737 ( .A0(n572), .A1(n571), .B0(n570), .Y(n573) );
  AO22X1 U738 ( .A0(\intadd_2/SUM[2] ), .A1(n539), .B0(IM_D[1]), .B1(n727), 
        .Y(n578) );
  AO22X1 U739 ( .A0(\intadd_2/SUM[3] ), .A1(n539), .B0(IM_D[2]), .B1(n727), 
        .Y(n581) );
  AO22X1 U740 ( .A0(\intadd_2/SUM[4] ), .A1(n539), .B0(IM_D[3]), .B1(n727), 
        .Y(n584) );
  AO22X1 U741 ( .A0(\intadd_2/SUM[5] ), .A1(n539), .B0(IM_D[4]), .B1(n727), 
        .Y(n587) );
  AO22X1 U742 ( .A0(\intadd_2/SUM[6] ), .A1(n539), .B0(IM_D[5]), .B1(n727), 
        .Y(n590) );
  OAI2BB2XL U743 ( .B0(n522), .B1(n466), .A0N(n640), .A1N(\intadd_2/SUM[5] ), 
        .Y(n593) );
  AOI2BB2X1 U744 ( .B0(im_d_w_9), .B1(n596), .A0N(im_d_w_9), .A1N(n596), .Y(
        n701) );
  OAI2BB2XL U745 ( .B0(n517), .B1(n466), .A0N(n640), .A1N(\intadd_2/SUM[6] ), 
        .Y(n597) );
  OAI21XL U746 ( .A0(\data_path/si_w[8] ), .A1(n615), .B0(en_so), .Y(n601) );
  AO22X1 U747 ( .A0(\intadd_1/SUM[6] ), .A1(n539), .B0(IM_D[13]), .B1(n727), 
        .Y(n605) );
  OAI2BB2XL U748 ( .B0(n466), .B1(n527), .A0N(n640), .A1N(\intadd_1/SUM[5] ), 
        .Y(n608) );
  AOI2BB2X1 U749 ( .B0(im_d_w_19), .B1(n611), .A0N(im_d_w_19), .A1N(n611), .Y(
        n729) );
  OAI2BB2XL U750 ( .B0(n466), .B1(n523), .A0N(n640), .A1N(\intadd_1/SUM[6] ), 
        .Y(n612) );
  OAI21XL U751 ( .A0(\data_path/si_w[16] ), .A1(n615), .B0(en_so), .Y(n616) );
  AO22X1 U752 ( .A0(\intadd_0/SUM[3] ), .A1(n539), .B0(IM_D[18]), .B1(n727), 
        .Y(n620) );
  AO22X1 U753 ( .A0(\intadd_0/SUM[4] ), .A1(n539), .B0(n779), .B1(n727), .Y(
        n623) );
  AO22X1 U754 ( .A0(\intadd_0/SUM[5] ), .A1(n539), .B0(n778), .B1(n727), .Y(
        n626) );
  AO22X1 U755 ( .A0(\intadd_0/SUM[6] ), .A1(n539), .B0(n777), .B1(n727), .Y(
        n630) );
  OAI2BB2XL U756 ( .B0(n466), .B1(n512), .A0N(n640), .A1N(\intadd_0/SUM[5] ), 
        .Y(n633) );
  AOI2BB2X1 U757 ( .B0(im_d_w[29]), .B1(n638), .A0N(im_d_w[29]), .A1N(n638), 
        .Y(n694) );
  OAI2BB2XL U758 ( .B0(n466), .B1(n513), .A0N(n640), .A1N(\intadd_0/SUM[6] ), 
        .Y(n642) );
  OAI22XL U759 ( .A0(curr_time[0]), .A1(n648), .B0(n515), .B1(n670), .Y(n647)
         );
  OAI21XL U760 ( .A0(n722), .A1(n498), .B0(n647), .Y(n336) );
  OAI22XL U761 ( .A0(en_init_time), .A1(n649), .B0(n722), .B1(n504), .Y(n650)
         );
  OAI21XL U762 ( .A0(n722), .A1(n516), .B0(n656), .Y(n335) );
  AO22X1 U763 ( .A0(n724), .A1(\data_path/si_w[6] ), .B0(n670), .B1(
        curr_time[6]), .Y(n333) );
  AO22X1 U764 ( .A0(n724), .A1(\data_path/si_w[7] ), .B0(n670), .B1(
        curr_time[7]), .Y(n332) );
  OAI21XL U765 ( .A0(n722), .A1(n500), .B0(n671), .Y(n331) );
  AOI2BB2X1 U766 ( .B0(n724), .B1(\data_path/si_w[16] ), .A0N(curr_time[16]), 
        .A1N(n686), .Y(n677) );
  OAI21XL U767 ( .A0(n721), .A1(n506), .B0(n677), .Y(n323) );
  OAI22XL U768 ( .A0(curr_time[17]), .A1(n681), .B0(n679), .B1(n682), .Y(n680)
         );
  OAI21XL U769 ( .A0(n722), .A1(n525), .B0(n680), .Y(n322) );
  OAI21XL U770 ( .A0(n683), .A1(n682), .B0(curr_time[18]), .Y(n684) );
  OAI22XL U771 ( .A0(curr_time[19]), .A1(n690), .B0(n535), .B1(n691), .Y(n689)
         );
  OAI21XL U772 ( .A0(n722), .A1(n526), .B0(n689), .Y(n320) );
  OAI22XL U773 ( .A0(n721), .A1(n534), .B0(n722), .B1(n511), .Y(n318) );
  OAI22XL U774 ( .A0(n721), .A1(n531), .B0(n722), .B1(n512), .Y(n317) );
  OAI22XL U775 ( .A0(n721), .A1(n503), .B0(n722), .B1(n513), .Y(n316) );
  AOI2BB2X1 U776 ( .B0(\data_path/si_w[9] ), .B1(n724), .A0N(curr_time[9]), 
        .A1N(n706), .Y(n700) );
  OAI21XL U777 ( .A0(n703), .A1(n529), .B0(n700), .Y(n330) );
  AOI2BB2X1 U778 ( .B0(n465), .B1(n521), .A0N(n465), .A1N(curr_photo_addr[9]), 
        .Y(n400) );
  AOI2BB2X1 U779 ( .B0(n464), .B1(n521), .A0N(n464), .A1N(fb_addr[9]), .Y(n401) );
  OAI21XL U780 ( .A0(curr_time[9]), .A1(n714), .B0(n703), .Y(n704) );
  AOI2BB2X1 U781 ( .B0(n465), .B1(n499), .A0N(n465), .A1N(curr_photo_addr[10]), 
        .Y(n397) );
  AOI2BB2X1 U782 ( .B0(n464), .B1(n499), .A0N(n464), .A1N(fb_addr[10]), .Y(
        n398) );
  AOI2BB1X1 U783 ( .A0N(n709), .A1N(n714), .B0(n723), .Y(n713) );
  AOI2BB2X1 U784 ( .B0(\data_path/si_w[11] ), .B1(n724), .A0N(curr_time[11]), 
        .A1N(n719), .Y(n711) );
  AOI2BB2X1 U785 ( .B0(n465), .B1(n501), .A0N(n465), .A1N(curr_photo_addr[11]), 
        .Y(n394) );
  AOI2BB2X1 U786 ( .B0(n464), .B1(n501), .A0N(n464), .A1N(fb_addr[11]), .Y(
        n395) );
  OAI21XL U787 ( .A0(curr_time[11]), .A1(n714), .B0(n713), .Y(n715) );
  AOI2BB2X1 U788 ( .B0(n465), .B1(n520), .A0N(n465), .A1N(curr_photo_addr[12]), 
        .Y(n391) );
  AOI2BB2X1 U789 ( .B0(n464), .B1(n520), .A0N(n464), .A1N(fb_addr[12]), .Y(
        n392) );
  AOI2BB2X1 U790 ( .B0(n465), .B1(n507), .A0N(n465), .A1N(curr_photo_addr[13]), 
        .Y(n388) );
  AOI2BB2X1 U791 ( .B0(n464), .B1(n507), .A0N(n464), .A1N(fb_addr[13]), .Y(
        n389) );
  AO22X1 U792 ( .A0(\data_path/si_w[13] ), .A1(n731), .B0(n541), .B1(IM_Q[13]), 
        .Y(n390) );
  AO22X1 U793 ( .A0(n724), .A1(\data_path/si_w[14] ), .B0(n723), .B1(
        curr_time[14]), .Y(n325) );
  AOI2BB2X1 U794 ( .B0(n465), .B1(n527), .A0N(n465), .A1N(curr_photo_addr[14]), 
        .Y(n385) );
  AOI2BB2X1 U795 ( .B0(n464), .B1(n527), .A0N(n464), .A1N(fb_addr[14]), .Y(
        n386) );
  AO22X1 U796 ( .A0(\data_path/si_w[14] ), .A1(n731), .B0(n541), .B1(IM_Q[14]), 
        .Y(n387) );
  AO22X1 U797 ( .A0(n724), .A1(\data_path/si_w[15] ), .B0(n723), .B1(
        curr_time[15]), .Y(n324) );
  AOI2BB2X1 U798 ( .B0(n465), .B1(n523), .A0N(n465), .A1N(curr_photo_addr[15]), 
        .Y(n382) );
  AOI2BB2X1 U799 ( .B0(n464), .B1(n523), .A0N(n464), .A1N(fb_addr[15]), .Y(
        n383) );
  AO22X1 U800 ( .A0(\data_path/si_w[15] ), .A1(n731), .B0(n541), .B1(IM_Q[15]), 
        .Y(n384) );
  AOI2BB2X1 U801 ( .B0(n465), .B1(n525), .A0N(n465), .A1N(curr_photo_addr[17]), 
        .Y(n379) );
  AOI2BB2X1 U802 ( .B0(n464), .B1(n525), .A0N(n464), .A1N(fb_addr[17]), .Y(
        n380) );
  AO22X1 U803 ( .A0(\data_path/si_w[17] ), .A1(n731), .B0(n541), .B1(IM_Q[17]), 
        .Y(n381) );
  AOI2BB2X1 U804 ( .B0(n465), .B1(n524), .A0N(n465), .A1N(curr_photo_addr[18]), 
        .Y(n376) );
  AOI2BB2X1 U805 ( .B0(n464), .B1(n524), .A0N(n464), .A1N(fb_addr[18]), .Y(
        n377) );
  AO22X1 U806 ( .A0(\data_path/si_w[18] ), .A1(n731), .B0(n541), .B1(IM_Q[18]), 
        .Y(n378) );
  AOI2BB2X1 U807 ( .B0(n465), .B1(n526), .A0N(n465), .A1N(curr_photo_addr[19]), 
        .Y(n373) );
  AOI2BB2X1 U808 ( .B0(n464), .B1(n526), .A0N(n464), .A1N(fb_addr[19]), .Y(
        n374) );
  AO22X1 U809 ( .A0(\data_path/si_w[19] ), .A1(n731), .B0(n541), .B1(IM_Q[19]), 
        .Y(n375) );
  AO22X1 U810 ( .A0(\data_path/si_w[20] ), .A1(n731), .B0(n541), .B1(IM_Q[20]), 
        .Y(n372) );
  AO22X1 U811 ( .A0(\data_path/si_w[21] ), .A1(n731), .B0(n541), .B1(IM_Q[21]), 
        .Y(n371) );
  AO22X1 U812 ( .A0(\data_path/si_w[22] ), .A1(n731), .B0(n541), .B1(IM_Q[22]), 
        .Y(n370) );
  AO22X1 U813 ( .A0(\data_path/si_w[23] ), .A1(n731), .B0(n541), .B1(IM_Q[23]), 
        .Y(n369) );
  AO22X1 U814 ( .A0(n465), .A1(\data_path/si_w[16] ), .B0(n543), .B1(
        curr_photo_addr[16]), .Y(n11) );
  AO22X1 U815 ( .A0(n464), .A1(\data_path/si_w[16] ), .B0(n544), .B1(
        fb_addr[16]), .Y(n12) );
  AOI2BB2X1 U816 ( .B0(n465), .B1(n500), .A0N(n465), .A1N(curr_photo_addr[8]), 
        .Y(n13) );
  AOI2BB2X1 U817 ( .B0(n464), .B1(n500), .A0N(n464), .A1N(fb_addr[8]), .Y(n14)
         );
  AOI2BB2X1 U818 ( .B0(n465), .B1(n509), .A0N(n465), .A1N(curr_photo_addr[4]), 
        .Y(n15) );
  AOI2BB2X1 U819 ( .B0(n464), .B1(n509), .A0N(n464), .A1N(fb_addr[4]), .Y(n16)
         );
  AOI2BB2X1 U820 ( .B0(n465), .B1(n510), .A0N(n465), .A1N(curr_photo_addr[2]), 
        .Y(n17) );
  AOI2BB2X1 U821 ( .B0(n464), .B1(n510), .A0N(n464), .A1N(fb_addr[2]), .Y(n18)
         );
  AOI2BB2X1 U822 ( .B0(n465), .B1(n504), .A0N(n465), .A1N(curr_photo_addr[1]), 
        .Y(n19) );
  AOI2BB2X1 U823 ( .B0(n464), .B1(n504), .A0N(n464), .A1N(fb_addr[1]), .Y(n20)
         );
  OAI22XL U824 ( .A0(\data_path/si_w[0] ), .A1(n504), .B0(n498), .B1(
        \data_path/si_w[1] ), .Y(n732) );
  OAI21XL U825 ( .A0(en_curr_photo_size), .A1(n530), .B0(n734), .Y(n23) );
endmodule

