
module p_dff_WORD20_NSEL5_0 ( clk, reset, en, sel, d, q );
  input [4:0] sel;
  input [19:0] d;
  output [19:0] q;
  input clk, reset, en;
  wire   n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31;

  DFFRX1 \q_reg[16]  ( .D(n60), .CK(clk), .RN(n31), .Q(q[16]) );
  DFFRX1 \q_reg[17]  ( .D(n61), .CK(clk), .RN(n31), .Q(q[17]) );
  DFFRX1 \q_reg[18]  ( .D(n62), .CK(clk), .RN(n31), .Q(q[18]) );
  DFFRX1 \q_reg[19]  ( .D(n63), .CK(clk), .RN(n31), .Q(q[19]) );
  DFFRX1 \q_reg[14]  ( .D(n58), .CK(clk), .RN(n31), .Q(q[14]) );
  DFFRX1 \q_reg[15]  ( .D(n59), .CK(clk), .RN(n31), .Q(q[15]) );
  DFFRX1 \q_reg[0]  ( .D(n44), .CK(clk), .RN(n31), .Q(q[0]) );
  DFFRX1 \q_reg[1]  ( .D(n45), .CK(clk), .RN(n31), .Q(q[1]) );
  DFFRX1 \q_reg[2]  ( .D(n46), .CK(clk), .RN(n31), .Q(q[2]) );
  DFFRX1 \q_reg[3]  ( .D(n47), .CK(clk), .RN(n31), .Q(q[3]) );
  DFFRX1 \q_reg[6]  ( .D(n50), .CK(clk), .RN(n31), .Q(q[6]) );
  DFFRX1 \q_reg[4]  ( .D(n48), .CK(clk), .RN(n31), .Q(q[4]) );
  DFFRX1 \q_reg[5]  ( .D(n49), .CK(clk), .RN(n31), .Q(q[5]) );
  DFFRX1 \q_reg[7]  ( .D(n51), .CK(clk), .RN(n31), .Q(q[7]) );
  DFFRX1 \q_reg[8]  ( .D(n52), .CK(clk), .RN(n31), .Q(q[8]) );
  DFFRX1 \q_reg[9]  ( .D(n53), .CK(clk), .RN(n31), .Q(q[9]) );
  DFFRX1 \q_reg[10]  ( .D(n54), .CK(clk), .RN(n31), .Q(q[10]) );
  DFFRX1 \q_reg[11]  ( .D(n55), .CK(clk), .RN(n31), .Q(q[11]) );
  DFFRX1 \q_reg[13]  ( .D(n57), .CK(clk), .RN(n31), .Q(q[13]) );
  DFFRX1 \q_reg[12]  ( .D(n56), .CK(clk), .RN(n31), .Q(q[12]) );
  INVX4 U3 ( .A(reset), .Y(n31) );
  INVX1 U4 ( .A(en), .Y(n6) );
  INVXL U5 ( .A(n13), .Y(n10) );
  MX2XL U6 ( .A(d[14]), .B(q[14]), .S0(n9), .Y(n58) );
  MX2X1 U7 ( .A(q[13]), .B(d[13]), .S0(n11), .Y(n57) );
  NOR2XL U8 ( .A(n8), .B(n9), .Y(n7) );
  MX2XL U9 ( .A(d[12]), .B(q[12]), .S0(n13), .Y(n56) );
  MX2XL U10 ( .A(q[4]), .B(d[4]), .S0(n25), .Y(n48) );
  MX2XL U11 ( .A(q[8]), .B(d[8]), .S0(n14), .Y(n52) );
  MX2XL U12 ( .A(d[6]), .B(q[6]), .S0(n24), .Y(n50) );
  CLKMX2X2 U13 ( .A(d[19]), .B(q[19]), .S0(n1), .Y(n63) );
  OAI31XL U14 ( .A0(sel[2]), .A1(sel[3]), .A2(sel[0]), .B0(n2), .Y(n1) );
  CLKMX2X2 U15 ( .A(q[18]), .B(d[18]), .S0(n2), .Y(n62) );
  OA21XL U16 ( .A0(sel[3]), .A1(n3), .B0(n4), .Y(n2) );
  CLKMX2X2 U17 ( .A(d[17]), .B(q[17]), .S0(n5), .Y(n61) );
  OAI31XL U18 ( .A0(sel[0]), .A1(sel[3]), .A2(n3), .B0(n4), .Y(n5) );
  CLKMX2X2 U19 ( .A(q[16]), .B(d[16]), .S0(n4), .Y(n60) );
  NOR2BX1 U20 ( .AN(sel[4]), .B(n6), .Y(n4) );
  CLKMX2X2 U21 ( .A(q[15]), .B(d[15]), .S0(n7), .Y(n59) );
  OAI21XL U22 ( .A0(sel[4]), .A1(sel[1]), .B0(n10), .Y(n9) );
  OA21XL U23 ( .A0(n12), .A1(sel[1]), .B0(n10), .Y(n11) );
  OAI21XL U24 ( .A0(sel[4]), .A1(sel[2]), .B0(n14), .Y(n13) );
  CLKMX2X2 U25 ( .A(q[11]), .B(d[11]), .S0(n15), .Y(n55) );
  AOI21X1 U26 ( .A0(n16), .A1(n17), .B0(n6), .Y(n15) );
  NAND3X1 U27 ( .A(sel[1]), .B(sel[0]), .C(sel[3]), .Y(n17) );
  OAI21XL U28 ( .A0(sel[4]), .A1(sel[2]), .B0(n18), .Y(n16) );
  CLKMX2X2 U29 ( .A(q[10]), .B(d[10]), .S0(n19), .Y(n54) );
  OA21XL U30 ( .A0(sel[4]), .A1(n3), .B0(n14), .Y(n19) );
  CLKMX2X2 U31 ( .A(q[9]), .B(d[9]), .S0(n20), .Y(n53) );
  OA21XL U32 ( .A0(n3), .A1(n12), .B0(n14), .Y(n20) );
  CLKINVX1 U33 ( .A(n8), .Y(n12) );
  NOR2X1 U34 ( .A(sel[0]), .B(sel[4]), .Y(n8) );
  NOR2X1 U35 ( .A(n6), .B(n21), .Y(n14) );
  CLKMX2X2 U36 ( .A(q[7]), .B(d[7]), .S0(n22), .Y(n51) );
  NOR2X1 U37 ( .A(n23), .B(n24), .Y(n22) );
  OAI21XL U38 ( .A0(sel[1]), .A1(n18), .B0(n25), .Y(n24) );
  CLKMX2X2 U39 ( .A(q[5]), .B(d[5]), .S0(n26), .Y(n49) );
  OA21XL U40 ( .A0(sel[1]), .A1(n27), .B0(n25), .Y(n26) );
  OA21XL U41 ( .A0(sel[2]), .A1(n18), .B0(en), .Y(n25) );
  CLKMX2X2 U42 ( .A(q[3]), .B(d[3]), .S0(n28), .Y(n47) );
  OA21XL U43 ( .A0(sel[2]), .A1(n27), .B0(n29), .Y(n28) );
  CLKMX2X2 U44 ( .A(q[2]), .B(d[2]), .S0(n29), .Y(n46) );
  OA21XL U45 ( .A0(n3), .A1(n18), .B0(en), .Y(n29) );
  CLKMX2X2 U46 ( .A(q[1]), .B(d[1]), .S0(n30), .Y(n45) );
  OA21XL U47 ( .A0(n3), .A1(n27), .B0(en), .Y(n30) );
  CLKINVX1 U48 ( .A(n23), .Y(n27) );
  NOR2X1 U49 ( .A(n18), .B(sel[0]), .Y(n23) );
  CLKINVX1 U50 ( .A(n21), .Y(n18) );
  NOR2X1 U51 ( .A(sel[3]), .B(sel[4]), .Y(n21) );
  OR2X1 U52 ( .A(sel[1]), .B(sel[2]), .Y(n3) );
  CLKMX2X2 U53 ( .A(d[0]), .B(q[0]), .S0(n6), .Y(n44) );
endmodule


module p_dff_WORD20_NSEL5_4 ( clk, reset, en, sel, d, q );
  input [4:0] sel;
  input [19:0] d;
  output [19:0] q;
  input clk, reset, en;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n52,
         n53, n54, n55, n56, n57, n58, n59;

  DFFRX1 \q_reg[19]  ( .D(n32), .CK(clk), .RN(n31), .Q(q[19]) );
  DFFRX1 \q_reg[17]  ( .D(n34), .CK(clk), .RN(n31), .Q(q[17]) );
  DFFRX1 \q_reg[18]  ( .D(n33), .CK(clk), .RN(n31), .Q(q[18]) );
  DFFRX1 \q_reg[16]  ( .D(n35), .CK(clk), .RN(n31), .Q(q[16]) );
  DFFRX1 \q_reg[15]  ( .D(n36), .CK(clk), .RN(n31), .Q(q[15]) );
  DFFRX1 \q_reg[14]  ( .D(n37), .CK(clk), .RN(n31), .Q(q[14]) );
  DFFRX1 \q_reg[12]  ( .D(n39), .CK(clk), .RN(n31), .Q(q[12]) );
  DFFRX1 \q_reg[13]  ( .D(n38), .CK(clk), .RN(n31), .Q(q[13]) );
  DFFRX1 \q_reg[11]  ( .D(n40), .CK(clk), .RN(n31), .Q(q[11]) );
  DFFRX1 \q_reg[10]  ( .D(n41), .CK(clk), .RN(n31), .Q(q[10]) );
  DFFRX1 \q_reg[9]  ( .D(n42), .CK(clk), .RN(n31), .Q(q[9]) );
  DFFRX1 \q_reg[6]  ( .D(n53), .CK(clk), .RN(n31), .Q(q[6]) );
  DFFRX1 \q_reg[8]  ( .D(n43), .CK(clk), .RN(n31), .Q(q[8]) );
  DFFRX1 \q_reg[7]  ( .D(n52), .CK(clk), .RN(n31), .Q(q[7]) );
  DFFRX1 \q_reg[5]  ( .D(n54), .CK(clk), .RN(n31), .Q(q[5]) );
  DFFRX1 \q_reg[4]  ( .D(n55), .CK(clk), .RN(n31), .Q(q[4]) );
  DFFRX1 \q_reg[3]  ( .D(n56), .CK(clk), .RN(n31), .Q(q[3]) );
  DFFRX1 \q_reg[2]  ( .D(n57), .CK(clk), .RN(n31), .Q(q[2]) );
  DFFRX2 \q_reg[0]  ( .D(n59), .CK(clk), .RN(n31), .Q(q[0]) );
  DFFRX2 \q_reg[1]  ( .D(n58), .CK(clk), .RN(n31), .Q(q[1]) );
  INVX4 U3 ( .A(reset), .Y(n31) );
  INVX1 U4 ( .A(en), .Y(n6) );
  INVXL U5 ( .A(n13), .Y(n10) );
  NOR2XL U6 ( .A(n8), .B(n9), .Y(n7) );
  MX2XL U7 ( .A(d[14]), .B(q[14]), .S0(n9), .Y(n37) );
  MX2XL U8 ( .A(d[12]), .B(q[12]), .S0(n13), .Y(n39) );
  MX2XL U9 ( .A(q[8]), .B(d[8]), .S0(n14), .Y(n43) );
  MX2XL U10 ( .A(d[6]), .B(q[6]), .S0(n24), .Y(n53) );
  NOR2XL U11 ( .A(n23), .B(n24), .Y(n22) );
  MX2XL U12 ( .A(q[4]), .B(d[4]), .S0(n25), .Y(n55) );
  CLKMX2X2 U13 ( .A(d[19]), .B(q[19]), .S0(n1), .Y(n32) );
  OAI31XL U14 ( .A0(sel[2]), .A1(sel[3]), .A2(sel[0]), .B0(n2), .Y(n1) );
  CLKMX2X2 U15 ( .A(q[18]), .B(d[18]), .S0(n2), .Y(n33) );
  OA21XL U16 ( .A0(sel[3]), .A1(n3), .B0(n4), .Y(n2) );
  CLKMX2X2 U17 ( .A(d[17]), .B(q[17]), .S0(n5), .Y(n34) );
  OAI31XL U18 ( .A0(sel[0]), .A1(sel[3]), .A2(n3), .B0(n4), .Y(n5) );
  CLKMX2X2 U19 ( .A(q[16]), .B(d[16]), .S0(n4), .Y(n35) );
  NOR2BX1 U20 ( .AN(sel[4]), .B(n6), .Y(n4) );
  CLKMX2X2 U21 ( .A(q[15]), .B(d[15]), .S0(n7), .Y(n36) );
  OAI21XL U22 ( .A0(sel[4]), .A1(sel[1]), .B0(n10), .Y(n9) );
  CLKMX2X2 U23 ( .A(q[13]), .B(d[13]), .S0(n11), .Y(n38) );
  OA21XL U24 ( .A0(n12), .A1(sel[1]), .B0(n10), .Y(n11) );
  OAI21XL U25 ( .A0(sel[4]), .A1(sel[2]), .B0(n14), .Y(n13) );
  CLKMX2X2 U26 ( .A(q[11]), .B(d[11]), .S0(n15), .Y(n40) );
  AOI21X1 U27 ( .A0(n16), .A1(n17), .B0(n6), .Y(n15) );
  NAND3X1 U28 ( .A(sel[1]), .B(sel[0]), .C(sel[3]), .Y(n17) );
  OAI21XL U29 ( .A0(sel[4]), .A1(sel[2]), .B0(n18), .Y(n16) );
  CLKMX2X2 U30 ( .A(q[10]), .B(d[10]), .S0(n19), .Y(n41) );
  OA21XL U31 ( .A0(sel[4]), .A1(n3), .B0(n14), .Y(n19) );
  CLKMX2X2 U32 ( .A(q[9]), .B(d[9]), .S0(n20), .Y(n42) );
  OA21XL U33 ( .A0(n3), .A1(n12), .B0(n14), .Y(n20) );
  CLKINVX1 U34 ( .A(n8), .Y(n12) );
  NOR2X1 U35 ( .A(sel[0]), .B(sel[4]), .Y(n8) );
  NOR2X1 U36 ( .A(n6), .B(n21), .Y(n14) );
  CLKMX2X2 U37 ( .A(q[7]), .B(d[7]), .S0(n22), .Y(n52) );
  OAI21XL U38 ( .A0(sel[1]), .A1(n18), .B0(n25), .Y(n24) );
  CLKMX2X2 U39 ( .A(q[5]), .B(d[5]), .S0(n26), .Y(n54) );
  OA21XL U40 ( .A0(sel[1]), .A1(n27), .B0(n25), .Y(n26) );
  OA21XL U41 ( .A0(sel[2]), .A1(n18), .B0(en), .Y(n25) );
  CLKMX2X2 U42 ( .A(q[3]), .B(d[3]), .S0(n28), .Y(n56) );
  OA21XL U43 ( .A0(sel[2]), .A1(n27), .B0(n29), .Y(n28) );
  CLKMX2X2 U44 ( .A(q[2]), .B(d[2]), .S0(n29), .Y(n57) );
  OA21XL U45 ( .A0(n3), .A1(n18), .B0(en), .Y(n29) );
  CLKMX2X2 U46 ( .A(q[1]), .B(d[1]), .S0(n30), .Y(n58) );
  OA21XL U47 ( .A0(n3), .A1(n27), .B0(en), .Y(n30) );
  CLKINVX1 U48 ( .A(n23), .Y(n27) );
  NOR2X1 U49 ( .A(n18), .B(sel[0]), .Y(n23) );
  CLKINVX1 U50 ( .A(n21), .Y(n18) );
  NOR2X1 U51 ( .A(sel[3]), .B(sel[4]), .Y(n21) );
  OR2X1 U52 ( .A(sel[1]), .B(sel[2]), .Y(n3) );
  CLKMX2X2 U53 ( .A(d[0]), .B(q[0]), .S0(n6), .Y(n59) );
endmodule


module p_dff_WORD9_NSEL4 ( clk, reset, en, sel, d, q );
  input [3:0] sel;
  input [8:0] d;
  output [8:0] q;
  input clk, reset, en;
  wire   n2, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n3, n4, n5, n6, n7, n8,
         n9, n32;

  DFFRHQX1 \q_reg[0]  ( .D(n23), .CK(clk), .RN(n32), .Q(q[0]) );
  DFFSRX1 \q_reg[5]  ( .D(n28), .CK(clk), .SN(1'b1), .RN(n32), .Q(q[5]), .QN(
        n2) );
  DFFRX1 \q_reg[8]  ( .D(n31), .CK(clk), .RN(n32), .Q(q[8]) );
  DFFRX1 \q_reg[4]  ( .D(n27), .CK(clk), .RN(n32), .Q(q[4]) );
  DFFRX1 \q_reg[6]  ( .D(n29), .CK(clk), .RN(n32), .Q(q[6]) );
  DFFRX1 \q_reg[2]  ( .D(n25), .CK(clk), .RN(n32), .Q(q[2]) );
  DFFRX1 \q_reg[1]  ( .D(n24), .CK(clk), .RN(n32), .Q(q[1]) );
  DFFRX1 \q_reg[7]  ( .D(n30), .CK(clk), .RN(n32), .Q(q[7]) );
  DFFRX1 \q_reg[3]  ( .D(n26), .CK(clk), .RN(n32), .Q(q[3]) );
  INVX1 U4 ( .A(en), .Y(n3) );
  CLKINVX1 U5 ( .A(n13), .Y(n5) );
  CLKINVX1 U6 ( .A(n20), .Y(n4) );
  INVX3 U7 ( .A(reset), .Y(n32) );
  OAI21X1 U8 ( .A0(sel[1]), .A1(n15), .B0(en), .Y(n13) );
  OAI21X1 U9 ( .A0(sel[3]), .A1(n19), .B0(en), .Y(n20) );
  NAND2X1 U10 ( .A(n10), .B(n11), .Y(n24) );
  NAND3BXL U11 ( .AN(n12), .B(en), .C(d[1]), .Y(n11) );
  OAI21XL U12 ( .A0(n12), .A1(n3), .B0(q[1]), .Y(n10) );
  NOR4X1 U13 ( .A(sel[0]), .B(sel[1]), .C(sel[2]), .D(sel[3]), .Y(n12) );
  OAI2BB2XL U14 ( .B0(n7), .B1(n16), .A0N(q[4]), .A1N(n16), .Y(n27) );
  CLKINVX1 U15 ( .A(d[4]), .Y(n7) );
  NAND2XL U16 ( .A(n15), .B(en), .Y(n16) );
  OAI2BB2XL U17 ( .B0(n9), .B1(n22), .A0N(q[8]), .A1N(n22), .Y(n31) );
  CLKINVX1 U18 ( .A(d[8]), .Y(n9) );
  NAND2XL U19 ( .A(sel[3]), .B(en), .Y(n22) );
  OAI2BB2XL U20 ( .B0(n6), .B1(n14), .A0N(q[3]), .A1N(n14), .Y(n26) );
  CLKINVX1 U21 ( .A(d[3]), .Y(n6) );
  OAI21X1 U22 ( .A0(sel[0]), .A1(n15), .B0(n5), .Y(n14) );
  OAI2BB2XL U23 ( .B0(n8), .B1(n21), .A0N(q[7]), .A1N(n21), .Y(n30) );
  CLKINVX1 U24 ( .A(d[7]), .Y(n8) );
  OAI21X1 U25 ( .A0(sel[3]), .A1(sel[0]), .B0(n4), .Y(n21) );
  OAI2BB2XL U26 ( .B0(n2), .B1(n17), .A0N(d[5]), .A1N(n17), .Y(n28) );
  NOR2X1 U27 ( .A(n18), .B(n3), .Y(n17) );
  AOI211X1 U28 ( .A0(sel[2]), .A1(sel[0]), .B0(n19), .C0(sel[3]), .Y(n18) );
  AO22XL U29 ( .A0(q[0]), .A1(n3), .B0(d[0]), .B1(en), .Y(n23) );
  AO22X1 U30 ( .A0(q[2]), .A1(n13), .B0(d[2]), .B1(n5), .Y(n25) );
  AO22X1 U31 ( .A0(q[6]), .A1(n20), .B0(d[6]), .B1(n4), .Y(n29) );
  OR2X1 U32 ( .A(sel[2]), .B(sel[3]), .Y(n15) );
  AND2X2 U33 ( .A(sel[1]), .B(sel[2]), .Y(n19) );
endmodule


module p_dff_WORD20_NSEL5_3 ( clk, reset, en, sel, d, q );
  input [4:0] sel;
  input [19:0] d;
  output [19:0] q;
  input clk, reset, en;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n52,
         n53, n54, n55, n56, n57, n58, n59;

  DFFRX1 \q_reg[2]  ( .D(n57), .CK(clk), .RN(n31), .Q(q[2]) );
  DFFRX1 \q_reg[1]  ( .D(n58), .CK(clk), .RN(n31), .Q(q[1]) );
  DFFRX1 \q_reg[0]  ( .D(n59), .CK(clk), .RN(n31), .Q(q[0]) );
  DFFRX1 \q_reg[5]  ( .D(n54), .CK(clk), .RN(n31), .Q(q[5]) );
  DFFRX1 \q_reg[4]  ( .D(n55), .CK(clk), .RN(n31), .Q(q[4]) );
  DFFRX1 \q_reg[3]  ( .D(n56), .CK(clk), .RN(n31), .Q(q[3]) );
  DFFRX2 \q_reg[14]  ( .D(n37), .CK(clk), .RN(n31), .Q(q[14]) );
  DFFRX2 \q_reg[17]  ( .D(n34), .CK(clk), .RN(n31), .Q(q[17]) );
  DFFRX2 \q_reg[18]  ( .D(n33), .CK(clk), .RN(n31), .Q(q[18]) );
  DFFRX2 \q_reg[19]  ( .D(n32), .CK(clk), .RN(n31), .Q(q[19]) );
  DFFRX2 \q_reg[16]  ( .D(n35), .CK(clk), .RN(n31), .Q(q[16]) );
  DFFRX2 \q_reg[7]  ( .D(n52), .CK(clk), .RN(n31), .Q(q[7]) );
  DFFRX2 \q_reg[15]  ( .D(n36), .CK(clk), .RN(n31), .Q(q[15]) );
  DFFRX2 \q_reg[10]  ( .D(n41), .CK(clk), .RN(n31), .Q(q[10]) );
  DFFRX2 \q_reg[13]  ( .D(n38), .CK(clk), .RN(n31), .Q(q[13]) );
  DFFRX2 \q_reg[11]  ( .D(n40), .CK(clk), .RN(n31), .Q(q[11]) );
  DFFRX2 \q_reg[6]  ( .D(n53), .CK(clk), .RN(n31), .Q(q[6]) );
  DFFRX2 \q_reg[8]  ( .D(n43), .CK(clk), .RN(n31), .Q(q[8]) );
  DFFRX2 \q_reg[9]  ( .D(n42), .CK(clk), .RN(n31), .Q(q[9]) );
  DFFRX2 \q_reg[12]  ( .D(n39), .CK(clk), .RN(n31), .Q(q[12]) );
  INVX4 U3 ( .A(reset), .Y(n31) );
  INVX1 U4 ( .A(en), .Y(n6) );
  INVXL U5 ( .A(n13), .Y(n10) );
  MX2XL U6 ( .A(d[14]), .B(q[14]), .S0(n9), .Y(n37) );
  MX2XL U7 ( .A(q[13]), .B(d[13]), .S0(n11), .Y(n38) );
  MX2XL U8 ( .A(q[9]), .B(d[9]), .S0(n20), .Y(n42) );
  MX2XL U9 ( .A(q[10]), .B(d[10]), .S0(n19), .Y(n41) );
  MX2XL U10 ( .A(d[12]), .B(q[12]), .S0(n13), .Y(n39) );
  MX2XL U11 ( .A(d[17]), .B(q[17]), .S0(n5), .Y(n34) );
  MX2XL U12 ( .A(q[18]), .B(d[18]), .S0(n2), .Y(n33) );
  MX2XL U13 ( .A(d[19]), .B(q[19]), .S0(n1), .Y(n32) );
  MX2XL U14 ( .A(q[16]), .B(d[16]), .S0(n4), .Y(n35) );
  MX2XL U15 ( .A(q[8]), .B(d[8]), .S0(n14), .Y(n43) );
  MX2XL U16 ( .A(q[11]), .B(d[11]), .S0(n15), .Y(n40) );
  MX2XL U17 ( .A(d[6]), .B(q[6]), .S0(n24), .Y(n53) );
  MX2XL U18 ( .A(q[4]), .B(d[4]), .S0(n25), .Y(n55) );
  MX2XL U19 ( .A(q[3]), .B(d[3]), .S0(n28), .Y(n56) );
  MX2XL U20 ( .A(q[5]), .B(d[5]), .S0(n26), .Y(n54) );
  MX2XL U21 ( .A(q[2]), .B(d[2]), .S0(n29), .Y(n57) );
  MX2XL U22 ( .A(q[1]), .B(d[1]), .S0(n30), .Y(n58) );
  MX2XL U23 ( .A(d[0]), .B(q[0]), .S0(n6), .Y(n59) );
  OAI31XL U24 ( .A0(sel[2]), .A1(sel[3]), .A2(sel[0]), .B0(n2), .Y(n1) );
  OA21XL U25 ( .A0(sel[3]), .A1(n3), .B0(n4), .Y(n2) );
  OAI31XL U26 ( .A0(sel[0]), .A1(sel[3]), .A2(n3), .B0(n4), .Y(n5) );
  NOR2BX1 U27 ( .AN(sel[4]), .B(n6), .Y(n4) );
  CLKMX2X2 U28 ( .A(q[15]), .B(d[15]), .S0(n7), .Y(n36) );
  NOR2X1 U29 ( .A(n8), .B(n9), .Y(n7) );
  OAI21XL U30 ( .A0(sel[4]), .A1(sel[1]), .B0(n10), .Y(n9) );
  OA21XL U31 ( .A0(n12), .A1(sel[1]), .B0(n10), .Y(n11) );
  OAI21XL U32 ( .A0(sel[4]), .A1(sel[2]), .B0(n14), .Y(n13) );
  AOI21X1 U33 ( .A0(n16), .A1(n17), .B0(n6), .Y(n15) );
  NAND3X1 U34 ( .A(sel[1]), .B(sel[0]), .C(sel[3]), .Y(n17) );
  OAI21XL U35 ( .A0(sel[4]), .A1(sel[2]), .B0(n18), .Y(n16) );
  OA21XL U36 ( .A0(sel[4]), .A1(n3), .B0(n14), .Y(n19) );
  OA21XL U37 ( .A0(n3), .A1(n12), .B0(n14), .Y(n20) );
  CLKINVX1 U38 ( .A(n8), .Y(n12) );
  NOR2X1 U39 ( .A(sel[0]), .B(sel[4]), .Y(n8) );
  NOR2X1 U40 ( .A(n6), .B(n21), .Y(n14) );
  CLKMX2X2 U41 ( .A(q[7]), .B(d[7]), .S0(n22), .Y(n52) );
  NOR2X1 U42 ( .A(n23), .B(n24), .Y(n22) );
  OAI21XL U43 ( .A0(sel[1]), .A1(n18), .B0(n25), .Y(n24) );
  OA21XL U44 ( .A0(sel[1]), .A1(n27), .B0(n25), .Y(n26) );
  OA21XL U45 ( .A0(sel[2]), .A1(n18), .B0(en), .Y(n25) );
  OA21XL U46 ( .A0(sel[2]), .A1(n27), .B0(n29), .Y(n28) );
  OA21XL U47 ( .A0(n3), .A1(n18), .B0(en), .Y(n29) );
  OA21XL U48 ( .A0(n3), .A1(n27), .B0(en), .Y(n30) );
  CLKINVX1 U49 ( .A(n23), .Y(n27) );
  NOR2X1 U50 ( .A(n18), .B(sel[0]), .Y(n23) );
  CLKINVX1 U51 ( .A(n21), .Y(n18) );
  NOR2X1 U52 ( .A(sel[3]), .B(sel[4]), .Y(n21) );
  OR2X1 U53 ( .A(sel[1]), .B(sel[2]), .Y(n3) );
endmodule


module CONT_DW_div_uns_0 ( a, b, quotient, remainder, divide_by_0 );
  input [19:0] a;
  input [3:0] b;
  output [19:0] quotient;
  output [3:0] remainder;
  output divide_by_0;
  wire   n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, \u_div/SumTmp[0][1] , \u_div/SumTmp[0][2] ,
         \u_div/SumTmp[0][3] , \u_div/SumTmp[1][1] , \u_div/SumTmp[1][2] ,
         \u_div/SumTmp[1][3] , \u_div/SumTmp[2][1] , \u_div/SumTmp[2][2] ,
         \u_div/SumTmp[2][3] , \u_div/SumTmp[3][1] , \u_div/SumTmp[3][2] ,
         \u_div/SumTmp[3][3] , \u_div/SumTmp[4][1] , \u_div/SumTmp[4][2] ,
         \u_div/SumTmp[4][3] , \u_div/SumTmp[5][1] , \u_div/SumTmp[5][2] ,
         \u_div/SumTmp[5][3] , \u_div/SumTmp[6][1] , \u_div/SumTmp[6][2] ,
         \u_div/SumTmp[6][3] , \u_div/SumTmp[7][1] , \u_div/SumTmp[7][2] ,
         \u_div/SumTmp[7][3] , \u_div/SumTmp[8][1] , \u_div/SumTmp[8][2] ,
         \u_div/SumTmp[8][3] , \u_div/SumTmp[9][1] , \u_div/SumTmp[9][2] ,
         \u_div/SumTmp[9][3] , \u_div/SumTmp[10][1] , \u_div/SumTmp[10][2] ,
         \u_div/SumTmp[10][3] , \u_div/SumTmp[11][1] , \u_div/SumTmp[11][2] ,
         \u_div/SumTmp[11][3] , \u_div/SumTmp[12][1] , \u_div/SumTmp[12][2] ,
         \u_div/SumTmp[12][3] , \u_div/SumTmp[13][1] , \u_div/SumTmp[13][2] ,
         \u_div/SumTmp[13][3] , \u_div/SumTmp[14][1] , \u_div/SumTmp[14][2] ,
         \u_div/SumTmp[14][3] , \u_div/SumTmp[15][1] , \u_div/SumTmp[15][2] ,
         \u_div/SumTmp[15][3] , \u_div/SumTmp[16][1] , \u_div/SumTmp[16][2] ,
         \u_div/SumTmp[16][3] , \u_div/CryTmp[0][1] , \u_div/CryTmp[1][1] ,
         \u_div/CryTmp[2][1] , \u_div/CryTmp[3][1] , \u_div/CryTmp[4][1] ,
         \u_div/CryTmp[5][1] , \u_div/CryTmp[6][1] , \u_div/CryTmp[7][1] ,
         \u_div/CryTmp[8][1] , \u_div/CryTmp[9][1] , \u_div/CryTmp[10][1] ,
         \u_div/CryTmp[11][1] , \u_div/CryTmp[12][1] , \u_div/CryTmp[13][1] ,
         \u_div/CryTmp[14][1] , \u_div/CryTmp[15][1] , \u_div/CryTmp[16][1] ,
         \u_div/CryTmp[17][1] , \u_div/CryTmp[18][1] , \u_div/PartRem[1][2] ,
         \u_div/PartRem[1][3] , \u_div/PartRem[2][1] , \u_div/PartRem[2][2] ,
         \u_div/PartRem[2][3] , \u_div/PartRem[3][1] , \u_div/PartRem[3][2] ,
         \u_div/PartRem[3][3] , \u_div/PartRem[4][1] , \u_div/PartRem[4][2] ,
         \u_div/PartRem[4][3] , \u_div/PartRem[5][1] , \u_div/PartRem[5][2] ,
         \u_div/PartRem[5][3] , \u_div/PartRem[6][1] , \u_div/PartRem[6][2] ,
         \u_div/PartRem[6][3] , \u_div/PartRem[7][1] , \u_div/PartRem[7][2] ,
         \u_div/PartRem[7][3] , \u_div/PartRem[8][1] , \u_div/PartRem[8][2] ,
         \u_div/PartRem[8][3] , \u_div/PartRem[9][1] , \u_div/PartRem[9][2] ,
         \u_div/PartRem[9][3] , \u_div/PartRem[10][1] , \u_div/PartRem[10][2] ,
         \u_div/PartRem[10][3] , \u_div/PartRem[11][1] ,
         \u_div/PartRem[11][2] , \u_div/PartRem[11][3] ,
         \u_div/PartRem[12][1] , \u_div/PartRem[12][2] ,
         \u_div/PartRem[12][3] , \u_div/PartRem[13][1] ,
         \u_div/PartRem[13][2] , \u_div/PartRem[13][3] ,
         \u_div/PartRem[14][1] , \u_div/PartRem[14][2] ,
         \u_div/PartRem[14][3] , \u_div/PartRem[15][1] ,
         \u_div/PartRem[15][2] , \u_div/PartRem[15][3] ,
         \u_div/PartRem[16][1] , \u_div/PartRem[16][2] ,
         \u_div/PartRem[16][3] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71;
  assign \u_div/CryTmp[0][1]  = a[0];
  assign \u_div/CryTmp[1][1]  = a[1];
  assign \u_div/CryTmp[2][1]  = a[2];
  assign \u_div/CryTmp[3][1]  = a[3];
  assign \u_div/CryTmp[4][1]  = a[4];
  assign \u_div/CryTmp[5][1]  = a[5];
  assign \u_div/CryTmp[6][1]  = a[6];
  assign \u_div/CryTmp[7][1]  = a[7];
  assign \u_div/CryTmp[8][1]  = a[8];
  assign \u_div/CryTmp[9][1]  = a[9];
  assign \u_div/CryTmp[10][1]  = a[10];
  assign \u_div/CryTmp[11][1]  = a[11];
  assign \u_div/CryTmp[12][1]  = a[12];
  assign \u_div/CryTmp[13][1]  = a[13];
  assign \u_div/CryTmp[14][1]  = a[14];
  assign \u_div/CryTmp[15][1]  = a[15];
  assign \u_div/CryTmp[16][1]  = a[16];
  assign \u_div/CryTmp[17][1]  = a[17];
  assign \u_div/CryTmp[18][1]  = a[18];

  MX2XL \u_div/u_mx_PartRem_0_0_1  ( .A(n2), .B(\u_div/SumTmp[0][1] ), .S0(n88), .Y(remainder[1]) );
  MX2X1 \u_div/u_mx_PartRem_0_16_2  ( .A(\u_div/CryTmp[18][1] ), .B(
        \u_div/SumTmp[16][2] ), .S0(n72), .Y(\u_div/PartRem[16][3] ) );
  MX2X1 \u_div/u_mx_PartRem_0_1_1  ( .A(\u_div/PartRem[2][1] ), .B(
        \u_div/SumTmp[1][1] ), .S0(n87), .Y(\u_div/PartRem[1][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_2_1  ( .A(\u_div/PartRem[3][1] ), .B(
        \u_div/SumTmp[2][1] ), .S0(n86), .Y(\u_div/PartRem[2][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_3_1  ( .A(\u_div/PartRem[4][1] ), .B(
        \u_div/SumTmp[3][1] ), .S0(n85), .Y(\u_div/PartRem[3][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_4_1  ( .A(\u_div/PartRem[5][1] ), .B(
        \u_div/SumTmp[4][1] ), .S0(n84), .Y(\u_div/PartRem[4][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_5_1  ( .A(\u_div/PartRem[6][1] ), .B(
        \u_div/SumTmp[5][1] ), .S0(n83), .Y(\u_div/PartRem[5][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_6_1  ( .A(\u_div/PartRem[7][1] ), .B(
        \u_div/SumTmp[6][1] ), .S0(n82), .Y(\u_div/PartRem[6][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_7_1  ( .A(\u_div/PartRem[8][1] ), .B(
        \u_div/SumTmp[7][1] ), .S0(n81), .Y(\u_div/PartRem[7][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_8_1  ( .A(\u_div/PartRem[9][1] ), .B(
        \u_div/SumTmp[8][1] ), .S0(n80), .Y(\u_div/PartRem[8][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_9_1  ( .A(\u_div/PartRem[10][1] ), .B(
        \u_div/SumTmp[9][1] ), .S0(n79), .Y(\u_div/PartRem[9][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_10_1  ( .A(\u_div/PartRem[11][1] ), .B(
        \u_div/SumTmp[10][1] ), .S0(n78), .Y(\u_div/PartRem[10][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_11_1  ( .A(\u_div/PartRem[12][1] ), .B(
        \u_div/SumTmp[11][1] ), .S0(n77), .Y(\u_div/PartRem[11][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_12_1  ( .A(\u_div/PartRem[13][1] ), .B(
        \u_div/SumTmp[12][1] ), .S0(n76), .Y(\u_div/PartRem[12][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_13_1  ( .A(\u_div/PartRem[14][1] ), .B(
        \u_div/SumTmp[13][1] ), .S0(n75), .Y(\u_div/PartRem[13][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_14_1  ( .A(\u_div/PartRem[15][1] ), .B(
        \u_div/SumTmp[14][1] ), .S0(n74), .Y(\u_div/PartRem[14][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_15_1  ( .A(\u_div/PartRem[16][1] ), .B(
        \u_div/SumTmp[15][1] ), .S0(n73), .Y(\u_div/PartRem[15][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_16_1  ( .A(\u_div/CryTmp[17][1] ), .B(
        \u_div/SumTmp[16][1] ), .S0(n72), .Y(\u_div/PartRem[16][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_0_2  ( .A(\u_div/PartRem[1][2] ), .B(
        \u_div/SumTmp[0][2] ), .S0(n88), .Y(remainder[2]) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_1_2  ( .A(\u_div/PartRem[2][2] ), .B(
        \u_div/SumTmp[1][2] ), .S0(n87), .Y(\u_div/PartRem[1][3] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_2_2  ( .A(\u_div/PartRem[3][2] ), .B(
        \u_div/SumTmp[2][2] ), .S0(n86), .Y(\u_div/PartRem[2][3] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_3_2  ( .A(\u_div/PartRem[4][2] ), .B(
        \u_div/SumTmp[3][2] ), .S0(n85), .Y(\u_div/PartRem[3][3] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_4_2  ( .A(\u_div/PartRem[5][2] ), .B(
        \u_div/SumTmp[4][2] ), .S0(n84), .Y(\u_div/PartRem[4][3] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_5_2  ( .A(\u_div/PartRem[6][2] ), .B(
        \u_div/SumTmp[5][2] ), .S0(n83), .Y(\u_div/PartRem[5][3] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_6_2  ( .A(\u_div/PartRem[7][2] ), .B(
        \u_div/SumTmp[6][2] ), .S0(n82), .Y(\u_div/PartRem[6][3] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_7_2  ( .A(\u_div/PartRem[8][2] ), .B(
        \u_div/SumTmp[7][2] ), .S0(n81), .Y(\u_div/PartRem[7][3] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_8_2  ( .A(\u_div/PartRem[9][2] ), .B(
        \u_div/SumTmp[8][2] ), .S0(n80), .Y(\u_div/PartRem[8][3] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_9_2  ( .A(\u_div/PartRem[10][2] ), .B(
        \u_div/SumTmp[9][2] ), .S0(n79), .Y(\u_div/PartRem[9][3] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_10_2  ( .A(\u_div/PartRem[11][2] ), .B(
        \u_div/SumTmp[10][2] ), .S0(n78), .Y(\u_div/PartRem[10][3] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_11_2  ( .A(\u_div/PartRem[12][2] ), .B(
        \u_div/SumTmp[11][2] ), .S0(n77), .Y(\u_div/PartRem[11][3] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_12_2  ( .A(\u_div/PartRem[13][2] ), .B(
        \u_div/SumTmp[12][2] ), .S0(n76), .Y(\u_div/PartRem[12][3] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_13_2  ( .A(\u_div/PartRem[14][2] ), .B(
        \u_div/SumTmp[13][2] ), .S0(n75), .Y(\u_div/PartRem[13][3] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_14_2  ( .A(\u_div/PartRem[15][2] ), .B(
        \u_div/SumTmp[14][2] ), .S0(n74), .Y(\u_div/PartRem[14][3] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_15_2  ( .A(\u_div/PartRem[16][2] ), .B(
        \u_div/SumTmp[15][2] ), .S0(n73), .Y(\u_div/PartRem[15][3] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_0_3  ( .A(\u_div/PartRem[1][3] ), .B(
        \u_div/SumTmp[0][3] ), .S0(n88), .Y(remainder[3]) );
  AO21X1 U1 ( .A0(n41), .A1(\u_div/PartRem[2][3] ), .B0(n1), .Y(n87) );
  CLKMX2X2 U2 ( .A(\u_div/PartRem[3][3] ), .B(\u_div/SumTmp[2][3] ), .S0(n86), 
        .Y(n1) );
  OR2X1 U3 ( .A(n4), .B(n5), .Y(n2) );
  MXI2X2 U4 ( .A(n28), .B(\u_div/CryTmp[16][1] ), .S0(n72), .Y(
        \u_div/PartRem[16][1] ) );
  AND2X2 U5 ( .A(a[19]), .B(n71), .Y(n72) );
  MXI2X2 U6 ( .A(n32), .B(\u_div/CryTmp[4][1] ), .S0(n84), .Y(
        \u_div/PartRem[4][1] ) );
  MXI2X2 U7 ( .A(n24), .B(\u_div/CryTmp[12][1] ), .S0(n76), .Y(
        \u_div/PartRem[12][1] ) );
  MXI2X2 U8 ( .A(n37), .B(\u_div/CryTmp[9][1] ), .S0(n79), .Y(
        \u_div/PartRem[9][1] ) );
  MXI2X2 U9 ( .A(n25), .B(\u_div/CryTmp[13][1] ), .S0(n75), .Y(
        \u_div/PartRem[13][1] ) );
  MXI2X2 U10 ( .A(n30), .B(\u_div/CryTmp[2][1] ), .S0(n86), .Y(
        \u_div/PartRem[2][1] ) );
  MXI2X2 U11 ( .A(n35), .B(\u_div/CryTmp[7][1] ), .S0(n81), .Y(
        \u_div/PartRem[7][1] ) );
  MXI2X2 U12 ( .A(n22), .B(\u_div/CryTmp[10][1] ), .S0(n78), .Y(
        \u_div/PartRem[10][1] ) );
  XNOR2XL U13 ( .A(\u_div/PartRem[9][1] ), .B(\u_div/CryTmp[8][1] ), .Y(
        \u_div/SumTmp[8][1] ) );
  MXI2X2 U14 ( .A(n36), .B(\u_div/CryTmp[8][1] ), .S0(n80), .Y(
        \u_div/PartRem[8][1] ) );
  XNOR2XL U15 ( .A(\u_div/PartRem[12][1] ), .B(\u_div/CryTmp[11][1] ), .Y(
        \u_div/SumTmp[11][1] ) );
  MXI2X2 U16 ( .A(n23), .B(\u_div/CryTmp[11][1] ), .S0(n77), .Y(
        \u_div/PartRem[11][1] ) );
  XNOR2XL U17 ( .A(\u_div/PartRem[7][1] ), .B(\u_div/CryTmp[6][1] ), .Y(
        \u_div/SumTmp[6][1] ) );
  MXI2X2 U18 ( .A(n34), .B(\u_div/CryTmp[6][1] ), .S0(n82), .Y(
        \u_div/PartRem[6][1] ) );
  XNOR2XL U19 ( .A(\u_div/PartRem[6][1] ), .B(\u_div/CryTmp[5][1] ), .Y(
        \u_div/SumTmp[5][1] ) );
  MXI2X2 U20 ( .A(n33), .B(\u_div/CryTmp[5][1] ), .S0(n83), .Y(
        \u_div/PartRem[5][1] ) );
  XNOR2XL U21 ( .A(\u_div/PartRem[4][1] ), .B(\u_div/CryTmp[3][1] ), .Y(
        \u_div/SumTmp[3][1] ) );
  MXI2X2 U22 ( .A(n31), .B(\u_div/CryTmp[3][1] ), .S0(n85), .Y(
        \u_div/PartRem[3][1] ) );
  INVXL U23 ( .A(n87), .Y(n3) );
  NOR2XL U24 ( .A(\u_div/CryTmp[1][1] ), .B(n3), .Y(n4) );
  NOR2XL U25 ( .A(n87), .B(n29), .Y(n5) );
  XNOR2XL U26 ( .A(n2), .B(\u_div/CryTmp[0][1] ), .Y(\u_div/SumTmp[0][1] ) );
  MXI2X2 U27 ( .A(n26), .B(\u_div/CryTmp[14][1] ), .S0(n74), .Y(
        \u_div/PartRem[14][1] ) );
  XNOR2XL U28 ( .A(\u_div/PartRem[16][1] ), .B(\u_div/CryTmp[15][1] ), .Y(
        \u_div/SumTmp[15][1] ) );
  MXI2X2 U29 ( .A(n27), .B(\u_div/CryTmp[15][1] ), .S0(n73), .Y(
        \u_div/PartRem[15][1] ) );
  INVXL U30 ( .A(\u_div/CryTmp[16][1] ), .Y(n28) );
  MXI2XL U31 ( .A(a[19]), .B(\u_div/SumTmp[16][3] ), .S0(n72), .Y(n20) );
  INVXL U32 ( .A(\u_div/CryTmp[0][1] ), .Y(n21) );
  OAI2BB1X1 U33 ( .A0N(n65), .A1N(\u_div/PartRem[14][3] ), .B0(n6), .Y(n75) );
  MXI2X1 U34 ( .A(\u_div/PartRem[15][3] ), .B(\u_div/SumTmp[14][3] ), .S0(n74), 
        .Y(n6) );
  OAI2BB1X1 U35 ( .A0N(n63), .A1N(\u_div/PartRem[13][3] ), .B0(n7), .Y(n76) );
  MXI2X1 U36 ( .A(\u_div/PartRem[14][3] ), .B(\u_div/SumTmp[13][3] ), .S0(n75), 
        .Y(n7) );
  OAI2BB1X1 U37 ( .A0N(n61), .A1N(\u_div/PartRem[12][3] ), .B0(n8), .Y(n77) );
  MXI2X1 U38 ( .A(\u_div/PartRem[13][3] ), .B(\u_div/SumTmp[12][3] ), .S0(n76), 
        .Y(n8) );
  OAI2BB1X1 U39 ( .A0N(n59), .A1N(\u_div/PartRem[11][3] ), .B0(n9), .Y(n78) );
  MXI2X1 U40 ( .A(\u_div/PartRem[12][3] ), .B(\u_div/SumTmp[11][3] ), .S0(n77), 
        .Y(n9) );
  OAI2BB1X1 U41 ( .A0N(n57), .A1N(\u_div/PartRem[10][3] ), .B0(n10), .Y(n79)
         );
  MXI2X1 U42 ( .A(\u_div/PartRem[11][3] ), .B(\u_div/SumTmp[10][3] ), .S0(n78), 
        .Y(n10) );
  OAI2BB1X1 U43 ( .A0N(n55), .A1N(\u_div/PartRem[9][3] ), .B0(n11), .Y(n80) );
  MXI2X1 U44 ( .A(\u_div/PartRem[10][3] ), .B(\u_div/SumTmp[9][3] ), .S0(n79), 
        .Y(n11) );
  OAI2BB1X1 U45 ( .A0N(n53), .A1N(\u_div/PartRem[8][3] ), .B0(n12), .Y(n81) );
  MXI2X1 U46 ( .A(\u_div/PartRem[9][3] ), .B(\u_div/SumTmp[8][3] ), .S0(n80), 
        .Y(n12) );
  OAI2BB1X1 U47 ( .A0N(n51), .A1N(\u_div/PartRem[7][3] ), .B0(n13), .Y(n82) );
  MXI2X1 U48 ( .A(\u_div/PartRem[8][3] ), .B(\u_div/SumTmp[7][3] ), .S0(n81), 
        .Y(n13) );
  OAI2BB1X1 U49 ( .A0N(n49), .A1N(\u_div/PartRem[6][3] ), .B0(n14), .Y(n83) );
  MXI2X1 U50 ( .A(\u_div/PartRem[7][3] ), .B(\u_div/SumTmp[6][3] ), .S0(n82), 
        .Y(n14) );
  OAI2BB1X1 U51 ( .A0N(n47), .A1N(\u_div/PartRem[5][3] ), .B0(n15), .Y(n84) );
  MXI2X1 U52 ( .A(\u_div/PartRem[6][3] ), .B(\u_div/SumTmp[5][3] ), .S0(n83), 
        .Y(n15) );
  OAI2BB1X1 U53 ( .A0N(n45), .A1N(\u_div/PartRem[4][3] ), .B0(n16), .Y(n85) );
  MXI2X1 U54 ( .A(\u_div/PartRem[5][3] ), .B(\u_div/SumTmp[4][3] ), .S0(n84), 
        .Y(n16) );
  OAI2BB1X1 U55 ( .A0N(n43), .A1N(\u_div/PartRem[3][3] ), .B0(n17), .Y(n86) );
  MXI2X1 U56 ( .A(\u_div/PartRem[4][3] ), .B(\u_div/SumTmp[3][3] ), .S0(n85), 
        .Y(n17) );
  OAI2BB1X1 U57 ( .A0N(n39), .A1N(\u_div/PartRem[1][3] ), .B0(n18), .Y(n88) );
  MXI2X1 U58 ( .A(\u_div/PartRem[2][3] ), .B(\u_div/SumTmp[1][3] ), .S0(n87), 
        .Y(n18) );
  OAI2BB1X1 U59 ( .A0N(n67), .A1N(\u_div/PartRem[15][3] ), .B0(n19), .Y(n74)
         );
  MXI2X1 U60 ( .A(\u_div/PartRem[16][3] ), .B(\u_div/SumTmp[15][3] ), .S0(n73), 
        .Y(n19) );
  OAI2BB1X1 U61 ( .A0N(n69), .A1N(\u_div/PartRem[16][3] ), .B0(n20), .Y(n73)
         );
  CLKINVX1 U62 ( .A(\u_div/CryTmp[14][1] ), .Y(n26) );
  CLKINVX1 U63 ( .A(\u_div/CryTmp[5][1] ), .Y(n33) );
  CLKINVX1 U64 ( .A(\u_div/CryTmp[4][1] ), .Y(n32) );
  CLKINVX1 U65 ( .A(\u_div/CryTmp[3][1] ), .Y(n31) );
  CLKINVX1 U66 ( .A(\u_div/CryTmp[12][1] ), .Y(n24) );
  CLKINVX1 U67 ( .A(\u_div/CryTmp[6][1] ), .Y(n34) );
  CLKINVX1 U68 ( .A(\u_div/CryTmp[13][1] ), .Y(n25) );
  CLKINVX1 U69 ( .A(\u_div/CryTmp[11][1] ), .Y(n23) );
  CLKINVX1 U70 ( .A(\u_div/CryTmp[10][1] ), .Y(n22) );
  CLKINVX1 U71 ( .A(\u_div/CryTmp[9][1] ), .Y(n37) );
  CLKINVX1 U72 ( .A(\u_div/CryTmp[8][1] ), .Y(n36) );
  CLKINVX1 U73 ( .A(\u_div/CryTmp[7][1] ), .Y(n35) );
  CLKINVX1 U74 ( .A(\u_div/CryTmp[15][1] ), .Y(n27) );
  CLKINVX1 U75 ( .A(\u_div/CryTmp[2][1] ), .Y(n30) );
  CLKINVX1 U76 ( .A(\u_div/CryTmp[1][1] ), .Y(n29) );
  MXI2X1 U77 ( .A(n21), .B(\u_div/CryTmp[0][1] ), .S0(n88), .Y(remainder[0])
         );
  NOR2X1 U78 ( .A(\u_div/CryTmp[0][1] ), .B(n2), .Y(n38) );
  NOR2BX1 U79 ( .AN(\u_div/PartRem[1][2] ), .B(n38), .Y(n39) );
  XNOR2X1 U80 ( .A(\u_div/PartRem[1][2] ), .B(n38), .Y(\u_div/SumTmp[0][2] )
         );
  XOR2X1 U81 ( .A(\u_div/PartRem[1][3] ), .B(n39), .Y(\u_div/SumTmp[0][3] ) );
  NOR2X1 U82 ( .A(\u_div/CryTmp[1][1] ), .B(\u_div/PartRem[2][1] ), .Y(n40) );
  NOR2BX1 U83 ( .AN(\u_div/PartRem[2][2] ), .B(n40), .Y(n41) );
  XNOR2X1 U84 ( .A(\u_div/PartRem[2][1] ), .B(\u_div/CryTmp[1][1] ), .Y(
        \u_div/SumTmp[1][1] ) );
  XNOR2X1 U85 ( .A(\u_div/PartRem[2][2] ), .B(n40), .Y(\u_div/SumTmp[1][2] )
         );
  XOR2X1 U86 ( .A(\u_div/PartRem[2][3] ), .B(n41), .Y(\u_div/SumTmp[1][3] ) );
  NOR2X1 U87 ( .A(\u_div/CryTmp[2][1] ), .B(\u_div/PartRem[3][1] ), .Y(n42) );
  NOR2BX1 U88 ( .AN(\u_div/PartRem[3][2] ), .B(n42), .Y(n43) );
  XNOR2X1 U89 ( .A(\u_div/PartRem[3][1] ), .B(\u_div/CryTmp[2][1] ), .Y(
        \u_div/SumTmp[2][1] ) );
  XNOR2X1 U90 ( .A(\u_div/PartRem[3][2] ), .B(n42), .Y(\u_div/SumTmp[2][2] )
         );
  XOR2X1 U91 ( .A(\u_div/PartRem[3][3] ), .B(n43), .Y(\u_div/SumTmp[2][3] ) );
  NOR2X1 U92 ( .A(\u_div/CryTmp[3][1] ), .B(\u_div/PartRem[4][1] ), .Y(n44) );
  NOR2BX1 U93 ( .AN(\u_div/PartRem[4][2] ), .B(n44), .Y(n45) );
  XNOR2X1 U94 ( .A(\u_div/PartRem[4][2] ), .B(n44), .Y(\u_div/SumTmp[3][2] )
         );
  XOR2X1 U95 ( .A(\u_div/PartRem[4][3] ), .B(n45), .Y(\u_div/SumTmp[3][3] ) );
  NOR2X1 U96 ( .A(\u_div/CryTmp[4][1] ), .B(\u_div/PartRem[5][1] ), .Y(n46) );
  NOR2BX1 U97 ( .AN(\u_div/PartRem[5][2] ), .B(n46), .Y(n47) );
  XNOR2X1 U98 ( .A(\u_div/PartRem[5][1] ), .B(\u_div/CryTmp[4][1] ), .Y(
        \u_div/SumTmp[4][1] ) );
  XNOR2X1 U99 ( .A(\u_div/PartRem[5][2] ), .B(n46), .Y(\u_div/SumTmp[4][2] )
         );
  XOR2X1 U100 ( .A(\u_div/PartRem[5][3] ), .B(n47), .Y(\u_div/SumTmp[4][3] )
         );
  NOR2X1 U101 ( .A(\u_div/CryTmp[5][1] ), .B(\u_div/PartRem[6][1] ), .Y(n48)
         );
  NOR2BX1 U102 ( .AN(\u_div/PartRem[6][2] ), .B(n48), .Y(n49) );
  XNOR2X1 U103 ( .A(\u_div/PartRem[6][2] ), .B(n48), .Y(\u_div/SumTmp[5][2] )
         );
  XOR2X1 U104 ( .A(\u_div/PartRem[6][3] ), .B(n49), .Y(\u_div/SumTmp[5][3] )
         );
  NOR2X1 U105 ( .A(\u_div/CryTmp[6][1] ), .B(\u_div/PartRem[7][1] ), .Y(n50)
         );
  NOR2BX1 U106 ( .AN(\u_div/PartRem[7][2] ), .B(n50), .Y(n51) );
  XNOR2X1 U107 ( .A(\u_div/PartRem[7][2] ), .B(n50), .Y(\u_div/SumTmp[6][2] )
         );
  XOR2X1 U108 ( .A(\u_div/PartRem[7][3] ), .B(n51), .Y(\u_div/SumTmp[6][3] )
         );
  NOR2X1 U109 ( .A(\u_div/CryTmp[7][1] ), .B(\u_div/PartRem[8][1] ), .Y(n52)
         );
  NOR2BX1 U110 ( .AN(\u_div/PartRem[8][2] ), .B(n52), .Y(n53) );
  XNOR2X1 U111 ( .A(\u_div/PartRem[8][1] ), .B(\u_div/CryTmp[7][1] ), .Y(
        \u_div/SumTmp[7][1] ) );
  XNOR2X1 U112 ( .A(\u_div/PartRem[8][2] ), .B(n52), .Y(\u_div/SumTmp[7][2] )
         );
  XOR2X1 U113 ( .A(\u_div/PartRem[8][3] ), .B(n53), .Y(\u_div/SumTmp[7][3] )
         );
  NOR2X1 U114 ( .A(\u_div/CryTmp[8][1] ), .B(\u_div/PartRem[9][1] ), .Y(n54)
         );
  NOR2BX1 U115 ( .AN(\u_div/PartRem[9][2] ), .B(n54), .Y(n55) );
  XNOR2X1 U116 ( .A(\u_div/PartRem[9][2] ), .B(n54), .Y(\u_div/SumTmp[8][2] )
         );
  XOR2X1 U117 ( .A(\u_div/PartRem[9][3] ), .B(n55), .Y(\u_div/SumTmp[8][3] )
         );
  NOR2X1 U118 ( .A(\u_div/CryTmp[9][1] ), .B(\u_div/PartRem[10][1] ), .Y(n56)
         );
  NOR2BX1 U119 ( .AN(\u_div/PartRem[10][2] ), .B(n56), .Y(n57) );
  XNOR2X1 U120 ( .A(\u_div/PartRem[10][1] ), .B(\u_div/CryTmp[9][1] ), .Y(
        \u_div/SumTmp[9][1] ) );
  XNOR2X1 U121 ( .A(\u_div/PartRem[10][2] ), .B(n56), .Y(\u_div/SumTmp[9][2] )
         );
  XOR2X1 U122 ( .A(\u_div/PartRem[10][3] ), .B(n57), .Y(\u_div/SumTmp[9][3] )
         );
  NOR2X1 U123 ( .A(\u_div/CryTmp[10][1] ), .B(\u_div/PartRem[11][1] ), .Y(n58)
         );
  NOR2BX1 U124 ( .AN(\u_div/PartRem[11][2] ), .B(n58), .Y(n59) );
  XNOR2X1 U125 ( .A(\u_div/PartRem[11][1] ), .B(\u_div/CryTmp[10][1] ), .Y(
        \u_div/SumTmp[10][1] ) );
  XNOR2X1 U126 ( .A(\u_div/PartRem[11][2] ), .B(n58), .Y(\u_div/SumTmp[10][2] ) );
  XOR2X1 U127 ( .A(\u_div/PartRem[11][3] ), .B(n59), .Y(\u_div/SumTmp[10][3] )
         );
  NOR2X1 U128 ( .A(\u_div/CryTmp[11][1] ), .B(\u_div/PartRem[12][1] ), .Y(n60)
         );
  NOR2BX1 U129 ( .AN(\u_div/PartRem[12][2] ), .B(n60), .Y(n61) );
  XNOR2X1 U130 ( .A(\u_div/PartRem[12][2] ), .B(n60), .Y(\u_div/SumTmp[11][2] ) );
  XOR2X1 U131 ( .A(\u_div/PartRem[12][3] ), .B(n61), .Y(\u_div/SumTmp[11][3] )
         );
  NOR2X1 U132 ( .A(\u_div/CryTmp[12][1] ), .B(\u_div/PartRem[13][1] ), .Y(n62)
         );
  NOR2BX1 U133 ( .AN(\u_div/PartRem[13][2] ), .B(n62), .Y(n63) );
  XNOR2X1 U134 ( .A(\u_div/PartRem[13][1] ), .B(\u_div/CryTmp[12][1] ), .Y(
        \u_div/SumTmp[12][1] ) );
  XNOR2X1 U135 ( .A(\u_div/PartRem[13][2] ), .B(n62), .Y(\u_div/SumTmp[12][2] ) );
  XOR2X1 U136 ( .A(\u_div/PartRem[13][3] ), .B(n63), .Y(\u_div/SumTmp[12][3] )
         );
  NOR2X1 U137 ( .A(\u_div/CryTmp[13][1] ), .B(\u_div/PartRem[14][1] ), .Y(n64)
         );
  NOR2BX1 U138 ( .AN(\u_div/PartRem[14][2] ), .B(n64), .Y(n65) );
  XNOR2X1 U139 ( .A(\u_div/PartRem[14][1] ), .B(\u_div/CryTmp[13][1] ), .Y(
        \u_div/SumTmp[13][1] ) );
  XNOR2X1 U140 ( .A(\u_div/PartRem[14][2] ), .B(n64), .Y(\u_div/SumTmp[13][2] ) );
  XOR2X1 U141 ( .A(\u_div/PartRem[14][3] ), .B(n65), .Y(\u_div/SumTmp[13][3] )
         );
  NOR2X1 U142 ( .A(\u_div/CryTmp[14][1] ), .B(\u_div/PartRem[15][1] ), .Y(n66)
         );
  NOR2BX1 U143 ( .AN(\u_div/PartRem[15][2] ), .B(n66), .Y(n67) );
  XNOR2X1 U144 ( .A(\u_div/PartRem[15][1] ), .B(\u_div/CryTmp[14][1] ), .Y(
        \u_div/SumTmp[14][1] ) );
  XNOR2X1 U145 ( .A(\u_div/PartRem[15][2] ), .B(n66), .Y(\u_div/SumTmp[14][2] ) );
  XOR2X1 U146 ( .A(\u_div/PartRem[15][3] ), .B(n67), .Y(\u_div/SumTmp[14][3] )
         );
  NOR2X1 U147 ( .A(\u_div/CryTmp[15][1] ), .B(\u_div/PartRem[16][1] ), .Y(n68)
         );
  NOR2BX1 U148 ( .AN(\u_div/PartRem[16][2] ), .B(n68), .Y(n69) );
  XNOR2X1 U149 ( .A(\u_div/PartRem[16][2] ), .B(n68), .Y(\u_div/SumTmp[15][2] ) );
  XOR2X1 U150 ( .A(\u_div/PartRem[16][3] ), .B(n69), .Y(\u_div/SumTmp[15][3] )
         );
  NOR2X1 U151 ( .A(\u_div/CryTmp[16][1] ), .B(\u_div/CryTmp[17][1] ), .Y(n70)
         );
  NOR2BX1 U152 ( .AN(\u_div/CryTmp[18][1] ), .B(n70), .Y(n71) );
  XNOR2X1 U153 ( .A(\u_div/CryTmp[17][1] ), .B(\u_div/CryTmp[16][1] ), .Y(
        \u_div/SumTmp[16][1] ) );
  XNOR2X1 U154 ( .A(\u_div/CryTmp[18][1] ), .B(n70), .Y(\u_div/SumTmp[16][2] )
         );
  XOR2X1 U155 ( .A(a[19]), .B(n71), .Y(\u_div/SumTmp[16][3] ) );
endmodule


module CONT_DW01_inc_0 ( A, SUM );
  input [9:0] A;
  output [9:0] SUM;

  wire   [9:2] carry;

  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .Y(SUM[8]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module CONT_DW01_inc_1 ( A, SUM );
  input [20:0] A;
  output [20:0] SUM;

  wire   [20:2] carry;

  ADDHXL U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  ADDHXL U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  ADDHXL U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_18 ( .A(A[18]), .B(carry[18]), .CO(carry[19]), .S(SUM[18]) );
  ADDHXL U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  ADDHXL U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  ADDHXL U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  ADDHXL U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHXL U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHXL U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHXL U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1_1_19 ( .A(A[19]), .B(carry[19]), .Y(SUM[19]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module CONT_DW_div_uns_1 ( a, b, quotient, remainder, divide_by_0 );
  input [7:0] a;
  input [3:0] b;
  output [7:0] quotient;
  output [3:0] remainder;
  output divide_by_0;
  wire   n14, n15, n16, n17, n18, \u_div/SumTmp[0][0] , \u_div/SumTmp[0][2] ,
         \u_div/SumTmp[0][3] , \u_div/SumTmp[1][0] , \u_div/SumTmp[1][2] ,
         \u_div/SumTmp[1][3] , \u_div/SumTmp[2][0] , \u_div/SumTmp[2][2] ,
         \u_div/SumTmp[2][3] , \u_div/SumTmp[3][0] , \u_div/SumTmp[3][2] ,
         \u_div/SumTmp[3][3] , \u_div/SumTmp[4][0] , \u_div/SumTmp[4][2] ,
         \u_div/SumTmp[4][3] , \u_div/SumTmp[5][0] , \u_div/SumTmp[6][0] ,
         \u_div/SumTmp[7][0] , \u_div/PartRem[1][1] , \u_div/PartRem[1][2] ,
         \u_div/PartRem[1][3] , \u_div/PartRem[2][1] , \u_div/PartRem[2][2] ,
         \u_div/PartRem[2][3] , \u_div/PartRem[3][1] , \u_div/PartRem[3][2] ,
         \u_div/PartRem[3][3] , \u_div/PartRem[3][4] , \u_div/PartRem[4][1] ,
         \u_div/PartRem[4][2] , \u_div/PartRem[4][3] , n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13;
  assign \u_div/SumTmp[0][0]  = a[0];
  assign \u_div/SumTmp[1][0]  = a[1];
  assign \u_div/SumTmp[2][0]  = a[2];
  assign \u_div/SumTmp[3][0]  = a[3];
  assign \u_div/SumTmp[4][0]  = a[4];
  assign \u_div/SumTmp[5][0]  = a[5];
  assign \u_div/SumTmp[6][0]  = a[6];
  assign \u_div/SumTmp[7][0]  = a[7];

  MX2X1 \u_div/u_mx_PartRem_0_4_1  ( .A(\u_div/SumTmp[5][0] ), .B(n8), .S0(n14), .Y(\u_div/PartRem[4][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_4_2  ( .A(\u_div/SumTmp[6][0] ), .B(
        \u_div/SumTmp[4][2] ), .S0(n14), .Y(\u_div/PartRem[4][3] ) );
  MX2X1 \u_div/u_mx_PartRem_0_1_0  ( .A(\u_div/SumTmp[1][0] ), .B(
        \u_div/SumTmp[1][0] ), .S0(n17), .Y(\u_div/PartRem[1][1] ) );
  MX2X1 \u_div/u_mx_PartRem_0_2_0  ( .A(\u_div/SumTmp[2][0] ), .B(
        \u_div/SumTmp[2][0] ), .S0(n16), .Y(\u_div/PartRem[2][1] ) );
  MX2X1 \u_div/u_mx_PartRem_0_3_0  ( .A(\u_div/SumTmp[3][0] ), .B(
        \u_div/SumTmp[3][0] ), .S0(n15), .Y(\u_div/PartRem[3][1] ) );
  MX2X1 \u_div/u_mx_PartRem_0_0_0  ( .A(\u_div/SumTmp[0][0] ), .B(
        \u_div/SumTmp[0][0] ), .S0(n18), .Y(remainder[0]) );
  MX2X1 \u_div/u_mx_PartRem_0_4_0  ( .A(\u_div/SumTmp[4][0] ), .B(
        \u_div/SumTmp[4][0] ), .S0(n14), .Y(\u_div/PartRem[4][1] ) );
  MX2XL \u_div/u_mx_PartRem_0_0_1  ( .A(\u_div/PartRem[1][1] ), .B(n4), .S0(
        n18), .Y(remainder[1]) );
  MX2X1 \u_div/u_mx_PartRem_0_1_1  ( .A(\u_div/PartRem[2][1] ), .B(n5), .S0(
        n17), .Y(\u_div/PartRem[1][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_2_1  ( .A(\u_div/PartRem[3][1] ), .B(n6), .S0(
        n16), .Y(\u_div/PartRem[2][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_3_1  ( .A(\u_div/PartRem[4][1] ), .B(n7), .S0(
        n15), .Y(\u_div/PartRem[3][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_3_2  ( .A(\u_div/PartRem[4][2] ), .B(
        \u_div/SumTmp[3][2] ), .S0(n15), .Y(\u_div/PartRem[3][3] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_3_3  ( .A(\u_div/PartRem[4][3] ), .B(
        \u_div/SumTmp[3][3] ), .S0(n15), .Y(\u_div/PartRem[3][4] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_0_3  ( .A(\u_div/PartRem[1][3] ), .B(
        \u_div/SumTmp[0][3] ), .S0(n18), .Y(remainder[3]) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_0_2  ( .A(\u_div/PartRem[1][2] ), .B(
        \u_div/SumTmp[0][2] ), .S0(n18), .Y(remainder[2]) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_1_2  ( .A(\u_div/PartRem[2][2] ), .B(
        \u_div/SumTmp[1][2] ), .S0(n17), .Y(\u_div/PartRem[1][3] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_2_2  ( .A(\u_div/PartRem[3][2] ), .B(
        \u_div/SumTmp[2][2] ), .S0(n16), .Y(\u_div/PartRem[2][3] ) );
  NOR2X1 U1 ( .A(\u_div/SumTmp[6][0] ), .B(\u_div/SumTmp[5][0] ), .Y(n13) );
  XNOR2XL U2 ( .A(\u_div/SumTmp[7][0] ), .B(n13), .Y(\u_div/SumTmp[4][3] ) );
  XNOR2XL U3 ( .A(\u_div/SumTmp[5][0] ), .B(\u_div/SumTmp[6][0] ), .Y(
        \u_div/SumTmp[4][2] ) );
  NOR2BX2 U4 ( .AN(\u_div/SumTmp[7][0] ), .B(n13), .Y(n14) );
  MXI2XL U5 ( .A(\u_div/SumTmp[7][0] ), .B(\u_div/SumTmp[4][3] ), .S0(n14), 
        .Y(n3) );
  OAI2BB1X1 U6 ( .A0N(\u_div/PartRem[2][3] ), .A1N(n10), .B0(n1), .Y(n17) );
  MXI2X1 U7 ( .A(\u_div/PartRem[3][3] ), .B(\u_div/SumTmp[2][3] ), .S0(n16), 
        .Y(n1) );
  OAI2BB1X1 U8 ( .A0N(\u_div/PartRem[1][3] ), .A1N(n9), .B0(n2), .Y(n18) );
  MXI2X1 U9 ( .A(\u_div/PartRem[2][3] ), .B(\u_div/SumTmp[1][3] ), .S0(n17), 
        .Y(n2) );
  CLKINVX1 U10 ( .A(\u_div/PartRem[4][1] ), .Y(n7) );
  CLKINVX1 U11 ( .A(\u_div/PartRem[3][1] ), .Y(n6) );
  CLKINVX1 U12 ( .A(\u_div/PartRem[2][1] ), .Y(n5) );
  CLKINVX1 U13 ( .A(\u_div/PartRem[1][1] ), .Y(n4) );
  OAI2BB1X1 U14 ( .A0N(\u_div/PartRem[4][3] ), .A1N(n12), .B0(n3), .Y(n15) );
  CLKINVX1 U15 ( .A(\u_div/SumTmp[5][0] ), .Y(n8) );
  OR2X1 U16 ( .A(\u_div/PartRem[1][2] ), .B(\u_div/PartRem[1][1] ), .Y(n9) );
  XOR2X1 U17 ( .A(n4), .B(\u_div/PartRem[1][2] ), .Y(\u_div/SumTmp[0][2] ) );
  XOR2X1 U18 ( .A(\u_div/PartRem[1][3] ), .B(n9), .Y(\u_div/SumTmp[0][3] ) );
  OR2X1 U19 ( .A(\u_div/PartRem[2][2] ), .B(\u_div/PartRem[2][1] ), .Y(n10) );
  XOR2X1 U20 ( .A(n5), .B(\u_div/PartRem[2][2] ), .Y(\u_div/SumTmp[1][2] ) );
  XOR2X1 U21 ( .A(\u_div/PartRem[2][3] ), .B(n10), .Y(\u_div/SumTmp[1][3] ) );
  OR2X1 U22 ( .A(\u_div/PartRem[3][2] ), .B(\u_div/PartRem[3][1] ), .Y(n11) );
  AO21X1 U23 ( .A0(\u_div/PartRem[3][3] ), .A1(n11), .B0(\u_div/PartRem[3][4] ), .Y(n16) );
  XOR2X1 U24 ( .A(n6), .B(\u_div/PartRem[3][2] ), .Y(\u_div/SumTmp[2][2] ) );
  XOR2X1 U25 ( .A(\u_div/PartRem[3][3] ), .B(n11), .Y(\u_div/SumTmp[2][3] ) );
  OR2X1 U26 ( .A(\u_div/PartRem[4][2] ), .B(\u_div/PartRem[4][1] ), .Y(n12) );
  XOR2X1 U27 ( .A(n7), .B(\u_div/PartRem[4][2] ), .Y(\u_div/SumTmp[3][2] ) );
  XOR2X1 U28 ( .A(\u_div/PartRem[4][3] ), .B(n12), .Y(\u_div/SumTmp[3][3] ) );
endmodule


module CONT_DW_div_uns_2 ( a, b, quotient, remainder, divide_by_0 );
  input [7:0] a;
  input [3:0] b;
  output [7:0] quotient;
  output [3:0] remainder;
  output divide_by_0;
  wire   n14, \u_div/SumTmp[1][0] , \u_div/SumTmp[1][2] , \u_div/SumTmp[1][3] ,
         \u_div/SumTmp[2][0] , \u_div/SumTmp[2][2] , \u_div/SumTmp[2][3] ,
         \u_div/SumTmp[3][0] , \u_div/SumTmp[3][2] , \u_div/SumTmp[3][3] ,
         \u_div/SumTmp[4][0] , \u_div/SumTmp[4][2] , \u_div/SumTmp[4][3] ,
         \u_div/SumTmp[5][0] , \u_div/SumTmp[6][0] , \u_div/SumTmp[7][0] ,
         \u_div/PartRem[1][1] , \u_div/PartRem[1][2] , \u_div/PartRem[1][3] ,
         \u_div/PartRem[2][1] , \u_div/PartRem[2][2] , \u_div/PartRem[2][3] ,
         \u_div/PartRem[3][1] , \u_div/PartRem[3][2] , \u_div/PartRem[3][3] ,
         \u_div/PartRem[4][1] , \u_div/PartRem[4][2] , \u_div/PartRem[4][3] ,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13;
  assign \u_div/SumTmp[1][0]  = a[1];
  assign \u_div/SumTmp[2][0]  = a[2];
  assign \u_div/SumTmp[3][0]  = a[3];
  assign \u_div/SumTmp[4][0]  = a[4];
  assign \u_div/SumTmp[5][0]  = a[5];
  assign \u_div/SumTmp[6][0]  = a[6];
  assign \u_div/SumTmp[7][0]  = a[7];

  MX2XL \u_div/u_mx_PartRem_0_1_0  ( .A(\u_div/SumTmp[1][0] ), .B(
        \u_div/SumTmp[1][0] ), .S0(quotient[1]), .Y(\u_div/PartRem[1][1] ) );
  MX2X1 \u_div/u_mx_PartRem_0_4_1  ( .A(\u_div/SumTmp[5][0] ), .B(n8), .S0(n14), .Y(\u_div/PartRem[4][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_4_2  ( .A(\u_div/SumTmp[6][0] ), .B(
        \u_div/SumTmp[4][2] ), .S0(n14), .Y(\u_div/PartRem[4][3] ) );
  MX2X1 \u_div/u_mx_PartRem_0_3_0  ( .A(\u_div/SumTmp[3][0] ), .B(
        \u_div/SumTmp[3][0] ), .S0(quotient[3]), .Y(\u_div/PartRem[3][1] ) );
  MX2X1 \u_div/u_mx_PartRem_0_4_0  ( .A(\u_div/SumTmp[4][0] ), .B(
        \u_div/SumTmp[4][0] ), .S0(n14), .Y(\u_div/PartRem[4][1] ) );
  MX2XL \u_div/u_mx_PartRem_0_1_1  ( .A(\u_div/PartRem[2][1] ), .B(n5), .S0(
        quotient[1]), .Y(\u_div/PartRem[1][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_2_1  ( .A(\u_div/PartRem[3][1] ), .B(n6), .S0(
        quotient[2]), .Y(\u_div/PartRem[2][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_3_1  ( .A(\u_div/PartRem[4][1] ), .B(n7), .S0(
        quotient[3]), .Y(\u_div/PartRem[3][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_3_2  ( .A(\u_div/PartRem[4][2] ), .B(
        \u_div/SumTmp[3][2] ), .S0(quotient[3]), .Y(\u_div/PartRem[3][3] ) );
  MX2XL \u_div/u_mx_PartRem_0_1_2  ( .A(\u_div/PartRem[2][2] ), .B(
        \u_div/SumTmp[1][2] ), .S0(quotient[1]), .Y(\u_div/PartRem[1][3] ) );
  MX2X1 \u_div/u_mx_PartRem_0_2_2  ( .A(\u_div/PartRem[3][2] ), .B(
        \u_div/SumTmp[2][2] ), .S0(quotient[2]), .Y(\u_div/PartRem[2][3] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_2_0  ( .A(\u_div/SumTmp[2][0] ), .B(
        \u_div/SumTmp[2][0] ), .S0(quotient[2]), .Y(\u_div/PartRem[2][1] ) );
  NOR2X1 U1 ( .A(\u_div/SumTmp[6][0] ), .B(\u_div/SumTmp[5][0] ), .Y(n13) );
  XNOR2XL U2 ( .A(\u_div/SumTmp[7][0] ), .B(n13), .Y(\u_div/SumTmp[4][3] ) );
  OAI2BB1X2 U3 ( .A0N(\u_div/PartRem[2][3] ), .A1N(n10), .B0(n1), .Y(
        quotient[1]) );
  MXI2X1 U4 ( .A(\u_div/PartRem[3][3] ), .B(\u_div/SumTmp[2][3] ), .S0(
        quotient[2]), .Y(n1) );
  OAI2BB1X2 U5 ( .A0N(\u_div/PartRem[3][3] ), .A1N(n11), .B0(n2), .Y(
        quotient[2]) );
  MXI2X1 U6 ( .A(\u_div/PartRem[4][3] ), .B(\u_div/SumTmp[3][3] ), .S0(
        quotient[3]), .Y(n2) );
  OAI2BB1X2 U7 ( .A0N(\u_div/PartRem[4][3] ), .A1N(n12), .B0(n4), .Y(
        quotient[3]) );
  NOR2BX2 U8 ( .AN(\u_div/SumTmp[7][0] ), .B(n13), .Y(n14) );
  MXI2XL U9 ( .A(\u_div/PartRem[2][3] ), .B(\u_div/SumTmp[1][3] ), .S0(
        quotient[1]), .Y(n3) );
  MXI2XL U10 ( .A(\u_div/SumTmp[7][0] ), .B(\u_div/SumTmp[4][3] ), .S0(n14), 
        .Y(n4) );
  NAND2X1 U11 ( .A(n3), .B(n9), .Y(quotient[0]) );
  CLKINVX1 U12 ( .A(\u_div/PartRem[4][1] ), .Y(n7) );
  CLKINVX1 U13 ( .A(\u_div/PartRem[3][1] ), .Y(n6) );
  CLKINVX1 U14 ( .A(\u_div/PartRem[2][1] ), .Y(n5) );
  CLKINVX1 U15 ( .A(\u_div/SumTmp[5][0] ), .Y(n8) );
  OAI21XL U16 ( .A0(\u_div/PartRem[1][1] ), .A1(\u_div/PartRem[1][2] ), .B0(
        \u_div/PartRem[1][3] ), .Y(n9) );
  OR2X1 U17 ( .A(\u_div/PartRem[2][2] ), .B(\u_div/PartRem[2][1] ), .Y(n10) );
  XOR2X1 U18 ( .A(n5), .B(\u_div/PartRem[2][2] ), .Y(\u_div/SumTmp[1][2] ) );
  XOR2X1 U19 ( .A(\u_div/PartRem[2][3] ), .B(n10), .Y(\u_div/SumTmp[1][3] ) );
  OR2X1 U20 ( .A(\u_div/PartRem[3][2] ), .B(\u_div/PartRem[3][1] ), .Y(n11) );
  XOR2X1 U21 ( .A(n6), .B(\u_div/PartRem[3][2] ), .Y(\u_div/SumTmp[2][2] ) );
  XOR2X1 U22 ( .A(\u_div/PartRem[3][3] ), .B(n11), .Y(\u_div/SumTmp[2][3] ) );
  OR2X1 U23 ( .A(\u_div/PartRem[4][2] ), .B(\u_div/PartRem[4][1] ), .Y(n12) );
  XOR2X1 U24 ( .A(n7), .B(\u_div/PartRem[4][2] ), .Y(\u_div/SumTmp[3][2] ) );
  XOR2X1 U25 ( .A(\u_div/PartRem[4][3] ), .B(n12), .Y(\u_div/SumTmp[3][3] ) );
  XNOR2X1 U26 ( .A(\u_div/SumTmp[5][0] ), .B(\u_div/SumTmp[6][0] ), .Y(
        \u_div/SumTmp[4][2] ) );
endmodule


module CONT_DW_div_uns_3 ( a, b, quotient, remainder, divide_by_0 );
  input [7:0] a;
  input [3:0] b;
  output [7:0] quotient;
  output [3:0] remainder;
  output divide_by_0;
  wire   n14, n15, n16, n17, n18, \u_div/SumTmp[0][0] , \u_div/SumTmp[0][2] ,
         \u_div/SumTmp[0][3] , \u_div/SumTmp[1][0] , \u_div/SumTmp[1][2] ,
         \u_div/SumTmp[1][3] , \u_div/SumTmp[2][0] , \u_div/SumTmp[2][2] ,
         \u_div/SumTmp[2][3] , \u_div/SumTmp[3][0] , \u_div/SumTmp[3][2] ,
         \u_div/SumTmp[3][3] , \u_div/SumTmp[4][0] , \u_div/SumTmp[4][2] ,
         \u_div/SumTmp[4][3] , \u_div/SumTmp[5][0] , \u_div/SumTmp[6][0] ,
         \u_div/SumTmp[7][0] , \u_div/PartRem[1][1] , \u_div/PartRem[1][2] ,
         \u_div/PartRem[1][3] , \u_div/PartRem[2][1] , \u_div/PartRem[2][2] ,
         \u_div/PartRem[2][3] , \u_div/PartRem[3][1] , \u_div/PartRem[3][2] ,
         \u_div/PartRem[3][3] , \u_div/PartRem[3][4] , \u_div/PartRem[4][1] ,
         \u_div/PartRem[4][2] , \u_div/PartRem[4][3] , n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13;
  assign \u_div/SumTmp[0][0]  = a[0];
  assign \u_div/SumTmp[1][0]  = a[1];
  assign \u_div/SumTmp[2][0]  = a[2];
  assign \u_div/SumTmp[3][0]  = a[3];
  assign \u_div/SumTmp[4][0]  = a[4];
  assign \u_div/SumTmp[5][0]  = a[5];
  assign \u_div/SumTmp[6][0]  = a[6];
  assign \u_div/SumTmp[7][0]  = a[7];

  MX2X1 \u_div/u_mx_PartRem_0_4_1  ( .A(\u_div/SumTmp[5][0] ), .B(n8), .S0(n14), .Y(\u_div/PartRem[4][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_4_2  ( .A(\u_div/SumTmp[6][0] ), .B(
        \u_div/SumTmp[4][2] ), .S0(n14), .Y(\u_div/PartRem[4][3] ) );
  MX2X1 \u_div/u_mx_PartRem_0_1_0  ( .A(\u_div/SumTmp[1][0] ), .B(
        \u_div/SumTmp[1][0] ), .S0(n17), .Y(\u_div/PartRem[1][1] ) );
  MX2X1 \u_div/u_mx_PartRem_0_2_0  ( .A(\u_div/SumTmp[2][0] ), .B(
        \u_div/SumTmp[2][0] ), .S0(n16), .Y(\u_div/PartRem[2][1] ) );
  MX2X1 \u_div/u_mx_PartRem_0_3_0  ( .A(\u_div/SumTmp[3][0] ), .B(
        \u_div/SumTmp[3][0] ), .S0(n15), .Y(\u_div/PartRem[3][1] ) );
  MX2X1 \u_div/u_mx_PartRem_0_0_0  ( .A(\u_div/SumTmp[0][0] ), .B(
        \u_div/SumTmp[0][0] ), .S0(n18), .Y(remainder[0]) );
  MX2X1 \u_div/u_mx_PartRem_0_4_0  ( .A(\u_div/SumTmp[4][0] ), .B(
        \u_div/SumTmp[4][0] ), .S0(n14), .Y(\u_div/PartRem[4][1] ) );
  MX2XL \u_div/u_mx_PartRem_0_0_1  ( .A(\u_div/PartRem[1][1] ), .B(n4), .S0(
        n18), .Y(remainder[1]) );
  MX2X1 \u_div/u_mx_PartRem_0_1_1  ( .A(\u_div/PartRem[2][1] ), .B(n5), .S0(
        n17), .Y(\u_div/PartRem[1][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_2_1  ( .A(\u_div/PartRem[3][1] ), .B(n6), .S0(
        n16), .Y(\u_div/PartRem[2][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_3_1  ( .A(\u_div/PartRem[4][1] ), .B(n7), .S0(
        n15), .Y(\u_div/PartRem[3][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_3_2  ( .A(\u_div/PartRem[4][2] ), .B(
        \u_div/SumTmp[3][2] ), .S0(n15), .Y(\u_div/PartRem[3][3] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_3_3  ( .A(\u_div/PartRem[4][3] ), .B(
        \u_div/SumTmp[3][3] ), .S0(n15), .Y(\u_div/PartRem[3][4] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_0_3  ( .A(\u_div/PartRem[1][3] ), .B(
        \u_div/SumTmp[0][3] ), .S0(n18), .Y(remainder[3]) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_0_2  ( .A(\u_div/PartRem[1][2] ), .B(
        \u_div/SumTmp[0][2] ), .S0(n18), .Y(remainder[2]) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_1_2  ( .A(\u_div/PartRem[2][2] ), .B(
        \u_div/SumTmp[1][2] ), .S0(n17), .Y(\u_div/PartRem[1][3] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_2_2  ( .A(\u_div/PartRem[3][2] ), .B(
        \u_div/SumTmp[2][2] ), .S0(n16), .Y(\u_div/PartRem[2][3] ) );
  NOR2X1 U1 ( .A(\u_div/SumTmp[6][0] ), .B(\u_div/SumTmp[5][0] ), .Y(n13) );
  XNOR2XL U2 ( .A(\u_div/SumTmp[7][0] ), .B(n13), .Y(\u_div/SumTmp[4][3] ) );
  XNOR2XL U3 ( .A(\u_div/SumTmp[5][0] ), .B(\u_div/SumTmp[6][0] ), .Y(
        \u_div/SumTmp[4][2] ) );
  NOR2BX2 U4 ( .AN(\u_div/SumTmp[7][0] ), .B(n13), .Y(n14) );
  MXI2XL U5 ( .A(\u_div/SumTmp[7][0] ), .B(\u_div/SumTmp[4][3] ), .S0(n14), 
        .Y(n3) );
  OAI2BB1X1 U6 ( .A0N(\u_div/PartRem[2][3] ), .A1N(n10), .B0(n1), .Y(n17) );
  MXI2X1 U7 ( .A(\u_div/PartRem[3][3] ), .B(\u_div/SumTmp[2][3] ), .S0(n16), 
        .Y(n1) );
  OAI2BB1X1 U8 ( .A0N(\u_div/PartRem[1][3] ), .A1N(n9), .B0(n2), .Y(n18) );
  MXI2X1 U9 ( .A(\u_div/PartRem[2][3] ), .B(\u_div/SumTmp[1][3] ), .S0(n17), 
        .Y(n2) );
  CLKINVX1 U10 ( .A(\u_div/PartRem[4][1] ), .Y(n7) );
  CLKINVX1 U11 ( .A(\u_div/PartRem[3][1] ), .Y(n6) );
  CLKINVX1 U12 ( .A(\u_div/PartRem[2][1] ), .Y(n5) );
  CLKINVX1 U13 ( .A(\u_div/PartRem[1][1] ), .Y(n4) );
  OAI2BB1X1 U14 ( .A0N(\u_div/PartRem[4][3] ), .A1N(n12), .B0(n3), .Y(n15) );
  CLKINVX1 U15 ( .A(\u_div/SumTmp[5][0] ), .Y(n8) );
  OR2X1 U16 ( .A(\u_div/PartRem[1][2] ), .B(\u_div/PartRem[1][1] ), .Y(n9) );
  XOR2X1 U17 ( .A(n4), .B(\u_div/PartRem[1][2] ), .Y(\u_div/SumTmp[0][2] ) );
  XOR2X1 U18 ( .A(\u_div/PartRem[1][3] ), .B(n9), .Y(\u_div/SumTmp[0][3] ) );
  OR2X1 U19 ( .A(\u_div/PartRem[2][2] ), .B(\u_div/PartRem[2][1] ), .Y(n10) );
  XOR2X1 U20 ( .A(n5), .B(\u_div/PartRem[2][2] ), .Y(\u_div/SumTmp[1][2] ) );
  XOR2X1 U21 ( .A(\u_div/PartRem[2][3] ), .B(n10), .Y(\u_div/SumTmp[1][3] ) );
  OR2X1 U22 ( .A(\u_div/PartRem[3][2] ), .B(\u_div/PartRem[3][1] ), .Y(n11) );
  AO21X1 U23 ( .A0(\u_div/PartRem[3][3] ), .A1(n11), .B0(\u_div/PartRem[3][4] ), .Y(n16) );
  XOR2X1 U24 ( .A(n6), .B(\u_div/PartRem[3][2] ), .Y(\u_div/SumTmp[2][2] ) );
  XOR2X1 U25 ( .A(\u_div/PartRem[3][3] ), .B(n11), .Y(\u_div/SumTmp[2][3] ) );
  OR2X1 U26 ( .A(\u_div/PartRem[4][2] ), .B(\u_div/PartRem[4][1] ), .Y(n12) );
  XOR2X1 U27 ( .A(n7), .B(\u_div/PartRem[4][2] ), .Y(\u_div/SumTmp[3][2] ) );
  XOR2X1 U28 ( .A(\u_div/PartRem[4][3] ), .B(n12), .Y(\u_div/SumTmp[3][3] ) );
endmodule


module CONT_DW_div_uns_4 ( a, b, quotient, remainder, divide_by_0 );
  input [7:0] a;
  input [3:0] b;
  output [7:0] quotient;
  output [3:0] remainder;
  output divide_by_0;
  wire   n14, \u_div/SumTmp[1][0] , \u_div/SumTmp[1][2] , \u_div/SumTmp[1][3] ,
         \u_div/SumTmp[2][0] , \u_div/SumTmp[2][2] , \u_div/SumTmp[2][3] ,
         \u_div/SumTmp[3][0] , \u_div/SumTmp[3][2] , \u_div/SumTmp[3][3] ,
         \u_div/SumTmp[4][0] , \u_div/SumTmp[4][2] , \u_div/SumTmp[4][3] ,
         \u_div/SumTmp[5][0] , \u_div/SumTmp[6][0] , \u_div/SumTmp[7][0] ,
         \u_div/PartRem[1][1] , \u_div/PartRem[1][2] , \u_div/PartRem[1][3] ,
         \u_div/PartRem[2][1] , \u_div/PartRem[2][2] , \u_div/PartRem[2][3] ,
         \u_div/PartRem[3][1] , \u_div/PartRem[3][2] , \u_div/PartRem[3][3] ,
         \u_div/PartRem[4][1] , \u_div/PartRem[4][2] , \u_div/PartRem[4][3] ,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13;
  assign \u_div/SumTmp[1][0]  = a[1];
  assign \u_div/SumTmp[2][0]  = a[2];
  assign \u_div/SumTmp[3][0]  = a[3];
  assign \u_div/SumTmp[4][0]  = a[4];
  assign \u_div/SumTmp[5][0]  = a[5];
  assign \u_div/SumTmp[6][0]  = a[6];
  assign \u_div/SumTmp[7][0]  = a[7];

  MX2XL \u_div/u_mx_PartRem_0_1_0  ( .A(\u_div/SumTmp[1][0] ), .B(
        \u_div/SumTmp[1][0] ), .S0(quotient[1]), .Y(\u_div/PartRem[1][1] ) );
  MX2X1 \u_div/u_mx_PartRem_0_4_1  ( .A(\u_div/SumTmp[5][0] ), .B(n8), .S0(n14), .Y(\u_div/PartRem[4][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_4_2  ( .A(\u_div/SumTmp[6][0] ), .B(
        \u_div/SumTmp[4][2] ), .S0(n14), .Y(\u_div/PartRem[4][3] ) );
  MX2X1 \u_div/u_mx_PartRem_0_3_0  ( .A(\u_div/SumTmp[3][0] ), .B(
        \u_div/SumTmp[3][0] ), .S0(quotient[3]), .Y(\u_div/PartRem[3][1] ) );
  MX2X1 \u_div/u_mx_PartRem_0_4_0  ( .A(\u_div/SumTmp[4][0] ), .B(
        \u_div/SumTmp[4][0] ), .S0(n14), .Y(\u_div/PartRem[4][1] ) );
  MX2XL \u_div/u_mx_PartRem_0_1_1  ( .A(\u_div/PartRem[2][1] ), .B(n5), .S0(
        quotient[1]), .Y(\u_div/PartRem[1][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_2_1  ( .A(\u_div/PartRem[3][1] ), .B(n6), .S0(
        quotient[2]), .Y(\u_div/PartRem[2][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_3_1  ( .A(\u_div/PartRem[4][1] ), .B(n7), .S0(
        quotient[3]), .Y(\u_div/PartRem[3][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_3_2  ( .A(\u_div/PartRem[4][2] ), .B(
        \u_div/SumTmp[3][2] ), .S0(quotient[3]), .Y(\u_div/PartRem[3][3] ) );
  MX2XL \u_div/u_mx_PartRem_0_1_2  ( .A(\u_div/PartRem[2][2] ), .B(
        \u_div/SumTmp[1][2] ), .S0(quotient[1]), .Y(\u_div/PartRem[1][3] ) );
  MX2X1 \u_div/u_mx_PartRem_0_2_2  ( .A(\u_div/PartRem[3][2] ), .B(
        \u_div/SumTmp[2][2] ), .S0(quotient[2]), .Y(\u_div/PartRem[2][3] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_2_0  ( .A(\u_div/SumTmp[2][0] ), .B(
        \u_div/SumTmp[2][0] ), .S0(quotient[2]), .Y(\u_div/PartRem[2][1] ) );
  NOR2X1 U1 ( .A(\u_div/SumTmp[6][0] ), .B(\u_div/SumTmp[5][0] ), .Y(n13) );
  XNOR2XL U2 ( .A(\u_div/SumTmp[7][0] ), .B(n13), .Y(\u_div/SumTmp[4][3] ) );
  OAI2BB1X2 U3 ( .A0N(\u_div/PartRem[2][3] ), .A1N(n10), .B0(n1), .Y(
        quotient[1]) );
  MXI2X1 U4 ( .A(\u_div/PartRem[3][3] ), .B(\u_div/SumTmp[2][3] ), .S0(
        quotient[2]), .Y(n1) );
  OAI2BB1X2 U5 ( .A0N(\u_div/PartRem[3][3] ), .A1N(n11), .B0(n2), .Y(
        quotient[2]) );
  MXI2X1 U6 ( .A(\u_div/PartRem[4][3] ), .B(\u_div/SumTmp[3][3] ), .S0(
        quotient[3]), .Y(n2) );
  OAI2BB1X2 U7 ( .A0N(\u_div/PartRem[4][3] ), .A1N(n12), .B0(n4), .Y(
        quotient[3]) );
  NOR2BX2 U8 ( .AN(\u_div/SumTmp[7][0] ), .B(n13), .Y(n14) );
  MXI2XL U9 ( .A(\u_div/PartRem[2][3] ), .B(\u_div/SumTmp[1][3] ), .S0(
        quotient[1]), .Y(n3) );
  MXI2XL U10 ( .A(\u_div/SumTmp[7][0] ), .B(\u_div/SumTmp[4][3] ), .S0(n14), 
        .Y(n4) );
  NAND2X1 U11 ( .A(n3), .B(n9), .Y(quotient[0]) );
  CLKINVX1 U12 ( .A(\u_div/PartRem[4][1] ), .Y(n7) );
  CLKINVX1 U13 ( .A(\u_div/PartRem[3][1] ), .Y(n6) );
  CLKINVX1 U14 ( .A(\u_div/PartRem[2][1] ), .Y(n5) );
  CLKINVX1 U15 ( .A(\u_div/SumTmp[5][0] ), .Y(n8) );
  OAI21XL U16 ( .A0(\u_div/PartRem[1][1] ), .A1(\u_div/PartRem[1][2] ), .B0(
        \u_div/PartRem[1][3] ), .Y(n9) );
  OR2X1 U17 ( .A(\u_div/PartRem[2][2] ), .B(\u_div/PartRem[2][1] ), .Y(n10) );
  XOR2X1 U18 ( .A(n5), .B(\u_div/PartRem[2][2] ), .Y(\u_div/SumTmp[1][2] ) );
  XOR2X1 U19 ( .A(\u_div/PartRem[2][3] ), .B(n10), .Y(\u_div/SumTmp[1][3] ) );
  OR2X1 U20 ( .A(\u_div/PartRem[3][2] ), .B(\u_div/PartRem[3][1] ), .Y(n11) );
  XOR2X1 U21 ( .A(n6), .B(\u_div/PartRem[3][2] ), .Y(\u_div/SumTmp[2][2] ) );
  XOR2X1 U22 ( .A(\u_div/PartRem[3][3] ), .B(n11), .Y(\u_div/SumTmp[2][3] ) );
  OR2X1 U23 ( .A(\u_div/PartRem[4][2] ), .B(\u_div/PartRem[4][1] ), .Y(n12) );
  XOR2X1 U24 ( .A(n7), .B(\u_div/PartRem[4][2] ), .Y(\u_div/SumTmp[3][2] ) );
  XOR2X1 U25 ( .A(\u_div/PartRem[4][3] ), .B(n12), .Y(\u_div/SumTmp[3][3] ) );
  XNOR2X1 U26 ( .A(\u_div/SumTmp[5][0] ), .B(\u_div/SumTmp[6][0] ), .Y(
        \u_div/SumTmp[4][2] ) );
endmodule


module CONT_DW_div_uns_5 ( a, b, quotient, remainder, divide_by_0 );
  input [7:0] a;
  input [3:0] b;
  output [7:0] quotient;
  output [3:0] remainder;
  output divide_by_0;
  wire   n14, n15, n16, n17, n18, \u_div/SumTmp[0][0] , \u_div/SumTmp[0][2] ,
         \u_div/SumTmp[0][3] , \u_div/SumTmp[1][0] , \u_div/SumTmp[1][2] ,
         \u_div/SumTmp[1][3] , \u_div/SumTmp[2][0] , \u_div/SumTmp[2][2] ,
         \u_div/SumTmp[2][3] , \u_div/SumTmp[3][0] , \u_div/SumTmp[3][2] ,
         \u_div/SumTmp[3][3] , \u_div/SumTmp[4][0] , \u_div/SumTmp[4][2] ,
         \u_div/SumTmp[4][3] , \u_div/SumTmp[5][0] , \u_div/SumTmp[6][0] ,
         \u_div/SumTmp[7][0] , \u_div/PartRem[1][1] , \u_div/PartRem[1][2] ,
         \u_div/PartRem[1][3] , \u_div/PartRem[2][1] , \u_div/PartRem[2][2] ,
         \u_div/PartRem[2][3] , \u_div/PartRem[3][1] , \u_div/PartRem[3][2] ,
         \u_div/PartRem[3][3] , \u_div/PartRem[3][4] , \u_div/PartRem[4][1] ,
         \u_div/PartRem[4][2] , \u_div/PartRem[4][3] , n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13;
  assign \u_div/SumTmp[0][0]  = a[0];
  assign \u_div/SumTmp[1][0]  = a[1];
  assign \u_div/SumTmp[2][0]  = a[2];
  assign \u_div/SumTmp[3][0]  = a[3];
  assign \u_div/SumTmp[4][0]  = a[4];
  assign \u_div/SumTmp[5][0]  = a[5];
  assign \u_div/SumTmp[6][0]  = a[6];
  assign \u_div/SumTmp[7][0]  = a[7];

  MX2X1 \u_div/u_mx_PartRem_0_4_1  ( .A(\u_div/SumTmp[5][0] ), .B(n8), .S0(n14), .Y(\u_div/PartRem[4][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_4_2  ( .A(\u_div/SumTmp[6][0] ), .B(
        \u_div/SumTmp[4][2] ), .S0(n14), .Y(\u_div/PartRem[4][3] ) );
  MX2X1 \u_div/u_mx_PartRem_0_1_0  ( .A(\u_div/SumTmp[1][0] ), .B(
        \u_div/SumTmp[1][0] ), .S0(n17), .Y(\u_div/PartRem[1][1] ) );
  MX2X1 \u_div/u_mx_PartRem_0_2_0  ( .A(\u_div/SumTmp[2][0] ), .B(
        \u_div/SumTmp[2][0] ), .S0(n16), .Y(\u_div/PartRem[2][1] ) );
  MX2X1 \u_div/u_mx_PartRem_0_3_0  ( .A(\u_div/SumTmp[3][0] ), .B(
        \u_div/SumTmp[3][0] ), .S0(n15), .Y(\u_div/PartRem[3][1] ) );
  MX2X1 \u_div/u_mx_PartRem_0_0_0  ( .A(\u_div/SumTmp[0][0] ), .B(
        \u_div/SumTmp[0][0] ), .S0(n18), .Y(remainder[0]) );
  MX2X1 \u_div/u_mx_PartRem_0_4_0  ( .A(\u_div/SumTmp[4][0] ), .B(
        \u_div/SumTmp[4][0] ), .S0(n14), .Y(\u_div/PartRem[4][1] ) );
  MX2XL \u_div/u_mx_PartRem_0_0_1  ( .A(\u_div/PartRem[1][1] ), .B(n4), .S0(
        n18), .Y(remainder[1]) );
  MX2X1 \u_div/u_mx_PartRem_0_1_1  ( .A(\u_div/PartRem[2][1] ), .B(n5), .S0(
        n17), .Y(\u_div/PartRem[1][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_2_1  ( .A(\u_div/PartRem[3][1] ), .B(n6), .S0(
        n16), .Y(\u_div/PartRem[2][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_3_1  ( .A(\u_div/PartRem[4][1] ), .B(n7), .S0(
        n15), .Y(\u_div/PartRem[3][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_3_2  ( .A(\u_div/PartRem[4][2] ), .B(
        \u_div/SumTmp[3][2] ), .S0(n15), .Y(\u_div/PartRem[3][3] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_3_3  ( .A(\u_div/PartRem[4][3] ), .B(
        \u_div/SumTmp[3][3] ), .S0(n15), .Y(\u_div/PartRem[3][4] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_0_3  ( .A(\u_div/PartRem[1][3] ), .B(
        \u_div/SumTmp[0][3] ), .S0(n18), .Y(remainder[3]) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_0_2  ( .A(\u_div/PartRem[1][2] ), .B(
        \u_div/SumTmp[0][2] ), .S0(n18), .Y(remainder[2]) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_1_2  ( .A(\u_div/PartRem[2][2] ), .B(
        \u_div/SumTmp[1][2] ), .S0(n17), .Y(\u_div/PartRem[1][3] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_2_2  ( .A(\u_div/PartRem[3][2] ), .B(
        \u_div/SumTmp[2][2] ), .S0(n16), .Y(\u_div/PartRem[2][3] ) );
  NOR2BX2 U1 ( .AN(\u_div/SumTmp[7][0] ), .B(n13), .Y(n14) );
  MXI2XL U2 ( .A(\u_div/SumTmp[7][0] ), .B(\u_div/SumTmp[4][3] ), .S0(n14), 
        .Y(n3) );
  OAI2BB1X1 U3 ( .A0N(\u_div/PartRem[2][3] ), .A1N(n10), .B0(n1), .Y(n17) );
  MXI2X1 U4 ( .A(\u_div/PartRem[3][3] ), .B(\u_div/SumTmp[2][3] ), .S0(n16), 
        .Y(n1) );
  OAI2BB1X1 U5 ( .A0N(\u_div/PartRem[1][3] ), .A1N(n9), .B0(n2), .Y(n18) );
  MXI2X1 U6 ( .A(\u_div/PartRem[2][3] ), .B(\u_div/SumTmp[1][3] ), .S0(n17), 
        .Y(n2) );
  CLKINVX1 U7 ( .A(\u_div/PartRem[4][1] ), .Y(n7) );
  CLKINVX1 U8 ( .A(\u_div/PartRem[3][1] ), .Y(n6) );
  CLKINVX1 U9 ( .A(\u_div/PartRem[2][1] ), .Y(n5) );
  CLKINVX1 U10 ( .A(\u_div/PartRem[1][1] ), .Y(n4) );
  OAI2BB1X1 U11 ( .A0N(\u_div/PartRem[4][3] ), .A1N(n12), .B0(n3), .Y(n15) );
  CLKINVX1 U12 ( .A(\u_div/SumTmp[5][0] ), .Y(n8) );
  OR2X1 U13 ( .A(\u_div/PartRem[1][2] ), .B(\u_div/PartRem[1][1] ), .Y(n9) );
  XOR2X1 U14 ( .A(n4), .B(\u_div/PartRem[1][2] ), .Y(\u_div/SumTmp[0][2] ) );
  XOR2X1 U15 ( .A(\u_div/PartRem[1][3] ), .B(n9), .Y(\u_div/SumTmp[0][3] ) );
  OR2X1 U16 ( .A(\u_div/PartRem[2][2] ), .B(\u_div/PartRem[2][1] ), .Y(n10) );
  XOR2X1 U17 ( .A(n5), .B(\u_div/PartRem[2][2] ), .Y(\u_div/SumTmp[1][2] ) );
  XOR2X1 U18 ( .A(\u_div/PartRem[2][3] ), .B(n10), .Y(\u_div/SumTmp[1][3] ) );
  OR2X1 U19 ( .A(\u_div/PartRem[3][2] ), .B(\u_div/PartRem[3][1] ), .Y(n11) );
  AO21X1 U20 ( .A0(\u_div/PartRem[3][3] ), .A1(n11), .B0(\u_div/PartRem[3][4] ), .Y(n16) );
  XOR2X1 U21 ( .A(n6), .B(\u_div/PartRem[3][2] ), .Y(\u_div/SumTmp[2][2] ) );
  XOR2X1 U22 ( .A(\u_div/PartRem[3][3] ), .B(n11), .Y(\u_div/SumTmp[2][3] ) );
  OR2X1 U23 ( .A(\u_div/PartRem[4][2] ), .B(\u_div/PartRem[4][1] ), .Y(n12) );
  XOR2X1 U24 ( .A(n7), .B(\u_div/PartRem[4][2] ), .Y(\u_div/SumTmp[3][2] ) );
  XOR2X1 U25 ( .A(\u_div/PartRem[4][3] ), .B(n12), .Y(\u_div/SumTmp[3][3] ) );
  NOR2X1 U26 ( .A(\u_div/SumTmp[6][0] ), .B(\u_div/SumTmp[5][0] ), .Y(n13) );
  XNOR2X1 U27 ( .A(\u_div/SumTmp[5][0] ), .B(\u_div/SumTmp[6][0] ), .Y(
        \u_div/SumTmp[4][2] ) );
  XNOR2X1 U28 ( .A(\u_div/SumTmp[7][0] ), .B(n13), .Y(\u_div/SumTmp[4][3] ) );
endmodule


module CONT_DW_div_uns_6 ( a, b, quotient, remainder, divide_by_0 );
  input [7:0] a;
  input [3:0] b;
  output [7:0] quotient;
  output [3:0] remainder;
  output divide_by_0;
  wire   n14, \u_div/SumTmp[1][0] , \u_div/SumTmp[1][2] , \u_div/SumTmp[1][3] ,
         \u_div/SumTmp[2][0] , \u_div/SumTmp[2][2] , \u_div/SumTmp[2][3] ,
         \u_div/SumTmp[3][0] , \u_div/SumTmp[3][2] , \u_div/SumTmp[3][3] ,
         \u_div/SumTmp[4][0] , \u_div/SumTmp[4][2] , \u_div/SumTmp[4][3] ,
         \u_div/SumTmp[5][0] , \u_div/SumTmp[6][0] , \u_div/SumTmp[7][0] ,
         \u_div/PartRem[1][1] , \u_div/PartRem[1][2] , \u_div/PartRem[1][3] ,
         \u_div/PartRem[2][1] , \u_div/PartRem[2][2] , \u_div/PartRem[2][3] ,
         \u_div/PartRem[3][1] , \u_div/PartRem[3][2] , \u_div/PartRem[3][3] ,
         \u_div/PartRem[4][1] , \u_div/PartRem[4][2] , \u_div/PartRem[4][3] ,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13;
  assign \u_div/SumTmp[1][0]  = a[1];
  assign \u_div/SumTmp[2][0]  = a[2];
  assign \u_div/SumTmp[3][0]  = a[3];
  assign \u_div/SumTmp[4][0]  = a[4];
  assign \u_div/SumTmp[5][0]  = a[5];
  assign \u_div/SumTmp[6][0]  = a[6];
  assign \u_div/SumTmp[7][0]  = a[7];

  MX2XL \u_div/u_mx_PartRem_0_1_0  ( .A(\u_div/SumTmp[1][0] ), .B(
        \u_div/SumTmp[1][0] ), .S0(quotient[1]), .Y(\u_div/PartRem[1][1] ) );
  MX2X1 \u_div/u_mx_PartRem_0_4_1  ( .A(\u_div/SumTmp[5][0] ), .B(n8), .S0(n14), .Y(\u_div/PartRem[4][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_4_2  ( .A(\u_div/SumTmp[6][0] ), .B(
        \u_div/SumTmp[4][2] ), .S0(n14), .Y(\u_div/PartRem[4][3] ) );
  MX2X1 \u_div/u_mx_PartRem_0_3_0  ( .A(\u_div/SumTmp[3][0] ), .B(
        \u_div/SumTmp[3][0] ), .S0(quotient[3]), .Y(\u_div/PartRem[3][1] ) );
  MX2X1 \u_div/u_mx_PartRem_0_4_0  ( .A(\u_div/SumTmp[4][0] ), .B(
        \u_div/SumTmp[4][0] ), .S0(n14), .Y(\u_div/PartRem[4][1] ) );
  MX2XL \u_div/u_mx_PartRem_0_1_1  ( .A(\u_div/PartRem[2][1] ), .B(n5), .S0(
        quotient[1]), .Y(\u_div/PartRem[1][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_2_1  ( .A(\u_div/PartRem[3][1] ), .B(n6), .S0(
        quotient[2]), .Y(\u_div/PartRem[2][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_3_1  ( .A(\u_div/PartRem[4][1] ), .B(n7), .S0(
        quotient[3]), .Y(\u_div/PartRem[3][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_3_2  ( .A(\u_div/PartRem[4][2] ), .B(
        \u_div/SumTmp[3][2] ), .S0(quotient[3]), .Y(\u_div/PartRem[3][3] ) );
  MX2XL \u_div/u_mx_PartRem_0_1_2  ( .A(\u_div/PartRem[2][2] ), .B(
        \u_div/SumTmp[1][2] ), .S0(quotient[1]), .Y(\u_div/PartRem[1][3] ) );
  MX2X1 \u_div/u_mx_PartRem_0_2_2  ( .A(\u_div/PartRem[3][2] ), .B(
        \u_div/SumTmp[2][2] ), .S0(quotient[2]), .Y(\u_div/PartRem[2][3] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_2_0  ( .A(\u_div/SumTmp[2][0] ), .B(
        \u_div/SumTmp[2][0] ), .S0(quotient[2]), .Y(\u_div/PartRem[2][1] ) );
  OAI2BB1X2 U1 ( .A0N(\u_div/PartRem[2][3] ), .A1N(n10), .B0(n1), .Y(
        quotient[1]) );
  MXI2X1 U2 ( .A(\u_div/PartRem[3][3] ), .B(\u_div/SumTmp[2][3] ), .S0(
        quotient[2]), .Y(n1) );
  OAI2BB1X2 U3 ( .A0N(\u_div/PartRem[3][3] ), .A1N(n11), .B0(n2), .Y(
        quotient[2]) );
  MXI2X1 U4 ( .A(\u_div/PartRem[4][3] ), .B(\u_div/SumTmp[3][3] ), .S0(
        quotient[3]), .Y(n2) );
  OAI2BB1X2 U5 ( .A0N(\u_div/PartRem[4][3] ), .A1N(n12), .B0(n4), .Y(
        quotient[3]) );
  NOR2BX2 U6 ( .AN(\u_div/SumTmp[7][0] ), .B(n13), .Y(n14) );
  MXI2XL U7 ( .A(\u_div/PartRem[2][3] ), .B(\u_div/SumTmp[1][3] ), .S0(
        quotient[1]), .Y(n3) );
  MXI2XL U8 ( .A(\u_div/SumTmp[7][0] ), .B(\u_div/SumTmp[4][3] ), .S0(n14), 
        .Y(n4) );
  NAND2X1 U9 ( .A(n3), .B(n9), .Y(quotient[0]) );
  CLKINVX1 U10 ( .A(\u_div/PartRem[2][1] ), .Y(n5) );
  CLKINVX1 U11 ( .A(\u_div/PartRem[4][1] ), .Y(n7) );
  CLKINVX1 U12 ( .A(\u_div/PartRem[3][1] ), .Y(n6) );
  CLKINVX1 U13 ( .A(\u_div/SumTmp[5][0] ), .Y(n8) );
  OAI21XL U14 ( .A0(\u_div/PartRem[1][1] ), .A1(\u_div/PartRem[1][2] ), .B0(
        \u_div/PartRem[1][3] ), .Y(n9) );
  OR2X1 U15 ( .A(\u_div/PartRem[2][2] ), .B(\u_div/PartRem[2][1] ), .Y(n10) );
  XOR2X1 U16 ( .A(n5), .B(\u_div/PartRem[2][2] ), .Y(\u_div/SumTmp[1][2] ) );
  XOR2X1 U17 ( .A(\u_div/PartRem[2][3] ), .B(n10), .Y(\u_div/SumTmp[1][3] ) );
  OR2X1 U18 ( .A(\u_div/PartRem[3][2] ), .B(\u_div/PartRem[3][1] ), .Y(n11) );
  XOR2X1 U19 ( .A(n6), .B(\u_div/PartRem[3][2] ), .Y(\u_div/SumTmp[2][2] ) );
  XOR2X1 U20 ( .A(\u_div/PartRem[3][3] ), .B(n11), .Y(\u_div/SumTmp[2][3] ) );
  OR2X1 U21 ( .A(\u_div/PartRem[4][2] ), .B(\u_div/PartRem[4][1] ), .Y(n12) );
  XOR2X1 U22 ( .A(n7), .B(\u_div/PartRem[4][2] ), .Y(\u_div/SumTmp[3][2] ) );
  XOR2X1 U23 ( .A(\u_div/PartRem[4][3] ), .B(n12), .Y(\u_div/SumTmp[3][3] ) );
  NOR2X1 U24 ( .A(\u_div/SumTmp[6][0] ), .B(\u_div/SumTmp[5][0] ), .Y(n13) );
  XNOR2X1 U25 ( .A(\u_div/SumTmp[5][0] ), .B(\u_div/SumTmp[6][0] ), .Y(
        \u_div/SumTmp[4][2] ) );
  XNOR2X1 U26 ( .A(\u_div/SumTmp[7][0] ), .B(n13), .Y(\u_div/SumTmp[4][3] ) );
endmodule


module CONT_DW_div_uns_8 ( a, b, quotient, remainder, divide_by_0 );
  input [19:0] a;
  input [3:0] b;
  output [19:0] quotient;
  output [3:0] remainder;
  output divide_by_0;
  wire   \u_div/SumTmp[1][1] , \u_div/SumTmp[1][2] , \u_div/SumTmp[1][3] ,
         \u_div/SumTmp[2][1] , \u_div/SumTmp[2][2] , \u_div/SumTmp[2][3] ,
         \u_div/SumTmp[3][1] , \u_div/SumTmp[3][2] , \u_div/SumTmp[3][3] ,
         \u_div/SumTmp[4][1] , \u_div/SumTmp[4][2] , \u_div/SumTmp[4][3] ,
         \u_div/SumTmp[5][1] , \u_div/SumTmp[5][2] , \u_div/SumTmp[5][3] ,
         \u_div/SumTmp[6][1] , \u_div/SumTmp[6][2] , \u_div/SumTmp[6][3] ,
         \u_div/SumTmp[7][1] , \u_div/SumTmp[7][2] , \u_div/SumTmp[7][3] ,
         \u_div/SumTmp[8][1] , \u_div/SumTmp[8][2] , \u_div/SumTmp[8][3] ,
         \u_div/SumTmp[9][1] , \u_div/SumTmp[9][2] , \u_div/SumTmp[9][3] ,
         \u_div/SumTmp[10][1] , \u_div/SumTmp[10][2] , \u_div/SumTmp[10][3] ,
         \u_div/SumTmp[11][1] , \u_div/SumTmp[11][2] , \u_div/SumTmp[11][3] ,
         \u_div/SumTmp[12][1] , \u_div/SumTmp[12][2] , \u_div/SumTmp[12][3] ,
         \u_div/SumTmp[13][1] , \u_div/SumTmp[13][2] , \u_div/SumTmp[13][3] ,
         \u_div/SumTmp[14][1] , \u_div/SumTmp[14][2] , \u_div/SumTmp[14][3] ,
         \u_div/SumTmp[15][1] , \u_div/SumTmp[15][2] , \u_div/SumTmp[15][3] ,
         \u_div/SumTmp[16][1] , \u_div/SumTmp[16][2] , \u_div/SumTmp[16][3] ,
         \u_div/CryTmp[0][1] , \u_div/CryTmp[1][1] , \u_div/CryTmp[2][1] ,
         \u_div/CryTmp[3][1] , \u_div/CryTmp[4][1] , \u_div/CryTmp[5][1] ,
         \u_div/CryTmp[6][1] , \u_div/CryTmp[7][1] , \u_div/CryTmp[8][1] ,
         \u_div/CryTmp[9][1] , \u_div/CryTmp[10][1] , \u_div/CryTmp[11][1] ,
         \u_div/CryTmp[12][1] , \u_div/CryTmp[13][1] , \u_div/CryTmp[14][1] ,
         \u_div/CryTmp[15][1] , \u_div/CryTmp[16][1] , \u_div/CryTmp[17][1] ,
         \u_div/CryTmp[18][1] , \u_div/PartRem[1][1] , \u_div/PartRem[1][2] ,
         \u_div/PartRem[1][3] , \u_div/PartRem[2][1] , \u_div/PartRem[2][2] ,
         \u_div/PartRem[2][3] , \u_div/PartRem[3][1] , \u_div/PartRem[3][2] ,
         \u_div/PartRem[3][3] , \u_div/PartRem[4][1] , \u_div/PartRem[4][2] ,
         \u_div/PartRem[4][3] , \u_div/PartRem[5][1] , \u_div/PartRem[5][2] ,
         \u_div/PartRem[5][3] , \u_div/PartRem[6][1] , \u_div/PartRem[6][2] ,
         \u_div/PartRem[6][3] , \u_div/PartRem[7][1] , \u_div/PartRem[7][2] ,
         \u_div/PartRem[7][3] , \u_div/PartRem[8][1] , \u_div/PartRem[8][2] ,
         \u_div/PartRem[8][3] , \u_div/PartRem[9][1] , \u_div/PartRem[9][2] ,
         \u_div/PartRem[9][3] , \u_div/PartRem[10][1] , \u_div/PartRem[10][2] ,
         \u_div/PartRem[10][3] , \u_div/PartRem[11][1] ,
         \u_div/PartRem[11][2] , \u_div/PartRem[11][3] ,
         \u_div/PartRem[12][1] , \u_div/PartRem[12][2] ,
         \u_div/PartRem[12][3] , \u_div/PartRem[13][2] ,
         \u_div/PartRem[13][3] , \u_div/PartRem[14][2] ,
         \u_div/PartRem[14][3] , \u_div/PartRem[15][1] ,
         \u_div/PartRem[15][2] , \u_div/PartRem[15][3] ,
         \u_div/PartRem[16][2] , \u_div/PartRem[16][3] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77;
  assign \u_div/CryTmp[0][1]  = a[0];
  assign \u_div/CryTmp[1][1]  = a[1];
  assign \u_div/CryTmp[2][1]  = a[2];
  assign \u_div/CryTmp[3][1]  = a[3];
  assign \u_div/CryTmp[4][1]  = a[4];
  assign \u_div/CryTmp[5][1]  = a[5];
  assign \u_div/CryTmp[6][1]  = a[6];
  assign \u_div/CryTmp[7][1]  = a[7];
  assign \u_div/CryTmp[8][1]  = a[8];
  assign \u_div/CryTmp[9][1]  = a[9];
  assign \u_div/CryTmp[10][1]  = a[10];
  assign \u_div/CryTmp[11][1]  = a[11];
  assign \u_div/CryTmp[12][1]  = a[12];
  assign \u_div/CryTmp[13][1]  = a[13];
  assign \u_div/CryTmp[14][1]  = a[14];
  assign \u_div/CryTmp[15][1]  = a[15];
  assign \u_div/CryTmp[16][1]  = a[16];
  assign \u_div/CryTmp[17][1]  = a[17];
  assign \u_div/CryTmp[18][1]  = a[18];

  MX2XL \u_div/u_mx_PartRem_0_1_1  ( .A(\u_div/PartRem[2][1] ), .B(
        \u_div/SumTmp[1][1] ), .S0(quotient[1]), .Y(\u_div/PartRem[1][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_13_1  ( .A(n3), .B(\u_div/SumTmp[13][1] ), .S0(
        quotient[13]), .Y(\u_div/PartRem[13][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_14_1  ( .A(\u_div/PartRem[15][1] ), .B(
        \u_div/SumTmp[14][1] ), .S0(quotient[14]), .Y(\u_div/PartRem[14][2] )
         );
  MX2X1 \u_div/u_mx_PartRem_0_15_1  ( .A(n2), .B(\u_div/SumTmp[15][1] ), .S0(
        quotient[15]), .Y(\u_div/PartRem[15][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_16_1  ( .A(\u_div/CryTmp[17][1] ), .B(
        \u_div/SumTmp[16][1] ), .S0(quotient[16]), .Y(\u_div/PartRem[16][2] )
         );
  MX2X1 \u_div/u_mx_PartRem_0_3_1  ( .A(\u_div/PartRem[4][1] ), .B(
        \u_div/SumTmp[3][1] ), .S0(quotient[3]), .Y(\u_div/PartRem[3][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_4_1  ( .A(\u_div/PartRem[5][1] ), .B(
        \u_div/SumTmp[4][1] ), .S0(quotient[4]), .Y(\u_div/PartRem[4][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_5_1  ( .A(\u_div/PartRem[6][1] ), .B(
        \u_div/SumTmp[5][1] ), .S0(quotient[5]), .Y(\u_div/PartRem[5][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_6_1  ( .A(\u_div/PartRem[7][1] ), .B(
        \u_div/SumTmp[6][1] ), .S0(quotient[6]), .Y(\u_div/PartRem[6][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_7_1  ( .A(\u_div/PartRem[8][1] ), .B(
        \u_div/SumTmp[7][1] ), .S0(quotient[7]), .Y(\u_div/PartRem[7][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_8_1  ( .A(\u_div/PartRem[9][1] ), .B(
        \u_div/SumTmp[8][1] ), .S0(quotient[8]), .Y(\u_div/PartRem[8][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_9_1  ( .A(\u_div/PartRem[10][1] ), .B(
        \u_div/SumTmp[9][1] ), .S0(quotient[9]), .Y(\u_div/PartRem[9][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_10_1  ( .A(\u_div/PartRem[11][1] ), .B(
        \u_div/SumTmp[10][1] ), .S0(quotient[10]), .Y(\u_div/PartRem[10][2] )
         );
  MX2X1 \u_div/u_mx_PartRem_0_11_1  ( .A(\u_div/PartRem[12][1] ), .B(
        \u_div/SumTmp[11][1] ), .S0(quotient[11]), .Y(\u_div/PartRem[11][2] )
         );
  MX2X1 \u_div/u_mx_PartRem_0_12_1  ( .A(n1), .B(\u_div/SumTmp[12][1] ), .S0(
        quotient[12]), .Y(\u_div/PartRem[12][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_13_2  ( .A(\u_div/PartRem[14][2] ), .B(
        \u_div/SumTmp[13][2] ), .S0(quotient[13]), .Y(\u_div/PartRem[13][3] )
         );
  MX2X1 \u_div/u_mx_PartRem_0_14_2  ( .A(\u_div/PartRem[15][2] ), .B(
        \u_div/SumTmp[14][2] ), .S0(quotient[14]), .Y(\u_div/PartRem[14][3] )
         );
  MX2X1 \u_div/u_mx_PartRem_0_15_2  ( .A(\u_div/PartRem[16][2] ), .B(
        \u_div/SumTmp[15][2] ), .S0(quotient[15]), .Y(\u_div/PartRem[15][3] )
         );
  MX2X1 \u_div/u_mx_PartRem_0_2_2  ( .A(\u_div/PartRem[3][2] ), .B(
        \u_div/SumTmp[2][2] ), .S0(quotient[2]), .Y(\u_div/PartRem[2][3] ) );
  MX2X1 \u_div/u_mx_PartRem_0_3_2  ( .A(\u_div/PartRem[4][2] ), .B(
        \u_div/SumTmp[3][2] ), .S0(quotient[3]), .Y(\u_div/PartRem[3][3] ) );
  MX2X1 \u_div/u_mx_PartRem_0_4_2  ( .A(\u_div/PartRem[5][2] ), .B(
        \u_div/SumTmp[4][2] ), .S0(quotient[4]), .Y(\u_div/PartRem[4][3] ) );
  MX2X1 \u_div/u_mx_PartRem_0_5_2  ( .A(\u_div/PartRem[6][2] ), .B(
        \u_div/SumTmp[5][2] ), .S0(quotient[5]), .Y(\u_div/PartRem[5][3] ) );
  MX2X1 \u_div/u_mx_PartRem_0_6_2  ( .A(\u_div/PartRem[7][2] ), .B(
        \u_div/SumTmp[6][2] ), .S0(quotient[6]), .Y(\u_div/PartRem[6][3] ) );
  MX2X1 \u_div/u_mx_PartRem_0_7_2  ( .A(\u_div/PartRem[8][2] ), .B(
        \u_div/SumTmp[7][2] ), .S0(quotient[7]), .Y(\u_div/PartRem[7][3] ) );
  MX2X1 \u_div/u_mx_PartRem_0_8_2  ( .A(\u_div/PartRem[9][2] ), .B(
        \u_div/SumTmp[8][2] ), .S0(quotient[8]), .Y(\u_div/PartRem[8][3] ) );
  MX2X1 \u_div/u_mx_PartRem_0_9_2  ( .A(\u_div/PartRem[10][2] ), .B(
        \u_div/SumTmp[9][2] ), .S0(quotient[9]), .Y(\u_div/PartRem[9][3] ) );
  MX2X1 \u_div/u_mx_PartRem_0_10_2  ( .A(\u_div/PartRem[11][2] ), .B(
        \u_div/SumTmp[10][2] ), .S0(quotient[10]), .Y(\u_div/PartRem[10][3] )
         );
  MX2X1 \u_div/u_mx_PartRem_0_11_2  ( .A(\u_div/PartRem[12][2] ), .B(
        \u_div/SumTmp[11][2] ), .S0(quotient[11]), .Y(\u_div/PartRem[11][3] )
         );
  MX2X1 \u_div/u_mx_PartRem_0_12_2  ( .A(\u_div/PartRem[13][2] ), .B(
        \u_div/SumTmp[12][2] ), .S0(quotient[12]), .Y(\u_div/PartRem[12][3] )
         );
  MX2XL \u_div/u_mx_PartRem_0_1_2  ( .A(\u_div/PartRem[2][2] ), .B(
        \u_div/SumTmp[1][2] ), .S0(quotient[1]), .Y(\u_div/PartRem[1][3] ) );
  MX2XL \u_div/u_mx_PartRem_0_16_2  ( .A(\u_div/CryTmp[18][1] ), .B(
        \u_div/SumTmp[16][2] ), .S0(quotient[16]), .Y(\u_div/PartRem[16][3] )
         );
  CLKMX2X2 \u_div/u_mx_PartRem_0_2_1  ( .A(\u_div/PartRem[3][1] ), .B(
        \u_div/SumTmp[2][1] ), .S0(quotient[2]), .Y(\u_div/PartRem[2][2] ) );
  AND2X2 U1 ( .A(a[19]), .B(n77), .Y(quotient[16]) );
  OR2X1 U2 ( .A(n5), .B(n6), .Y(n1) );
  OR2X1 U3 ( .A(n8), .B(n9), .Y(n2) );
  OR2X1 U4 ( .A(n11), .B(n12), .Y(n3) );
  MXI2X2 U5 ( .A(n31), .B(\u_div/CryTmp[12][1] ), .S0(quotient[12]), .Y(
        \u_div/PartRem[12][1] ) );
  MXI2X2 U6 ( .A(n39), .B(\u_div/CryTmp[4][1] ), .S0(quotient[4]), .Y(
        \u_div/PartRem[4][1] ) );
  MXI2X2 U7 ( .A(n44), .B(\u_div/CryTmp[9][1] ), .S0(quotient[9]), .Y(
        \u_div/PartRem[9][1] ) );
  MXI2X2 U8 ( .A(n42), .B(\u_div/CryTmp[7][1] ), .S0(quotient[7]), .Y(
        \u_div/PartRem[7][1] ) );
  XOR2XL U9 ( .A(\u_div/PartRem[16][3] ), .B(n75), .Y(\u_div/SumTmp[15][3] )
         );
  MXI2X2 U10 ( .A(n34), .B(\u_div/CryTmp[15][1] ), .S0(quotient[15]), .Y(
        \u_div/PartRem[15][1] ) );
  OAI2BB1X2 U11 ( .A0N(n75), .A1N(\u_div/PartRem[16][3] ), .B0(n27), .Y(
        quotient[15]) );
  OAI2BB1X2 U12 ( .A0N(n47), .A1N(\u_div/PartRem[2][3] ), .B0(n24), .Y(
        quotient[1]) );
  MXI2X2 U13 ( .A(n40), .B(\u_div/CryTmp[5][1] ), .S0(quotient[5]), .Y(
        \u_div/PartRem[5][1] ) );
  OAI2BB1X2 U14 ( .A0N(n55), .A1N(\u_div/PartRem[6][3] ), .B0(n20), .Y(
        quotient[5]) );
  MXI2X2 U15 ( .A(n29), .B(\u_div/CryTmp[10][1] ), .S0(quotient[10]), .Y(
        \u_div/PartRem[10][1] ) );
  OAI2BB1X2 U16 ( .A0N(n65), .A1N(\u_div/PartRem[11][3] ), .B0(n15), .Y(
        quotient[10]) );
  MXI2X2 U17 ( .A(n41), .B(\u_div/CryTmp[6][1] ), .S0(quotient[6]), .Y(
        \u_div/PartRem[6][1] ) );
  OAI2BB1X2 U18 ( .A0N(n57), .A1N(\u_div/PartRem[7][3] ), .B0(n19), .Y(
        quotient[6]) );
  OAI2BB1X2 U19 ( .A0N(n59), .A1N(\u_div/PartRem[8][3] ), .B0(n18), .Y(
        quotient[7]) );
  MXI2X2 U20 ( .A(n37), .B(\u_div/CryTmp[2][1] ), .S0(quotient[2]), .Y(
        \u_div/PartRem[2][1] ) );
  OAI2BB1X2 U21 ( .A0N(n49), .A1N(\u_div/PartRem[3][3] ), .B0(n23), .Y(
        quotient[2]) );
  INVXL U22 ( .A(quotient[13]), .Y(n4) );
  NOR2XL U23 ( .A(\u_div/CryTmp[13][1] ), .B(n4), .Y(n5) );
  NOR2XL U24 ( .A(quotient[13]), .B(n32), .Y(n6) );
  XNOR2XL U25 ( .A(n1), .B(\u_div/CryTmp[12][1] ), .Y(\u_div/SumTmp[12][1] )
         );
  OAI2BB1X2 U26 ( .A0N(n71), .A1N(\u_div/PartRem[14][3] ), .B0(n25), .Y(
        quotient[13]) );
  INVXL U27 ( .A(quotient[16]), .Y(n7) );
  NOR2XL U28 ( .A(\u_div/CryTmp[16][1] ), .B(n7), .Y(n8) );
  NOR2XL U29 ( .A(quotient[16]), .B(n35), .Y(n9) );
  XNOR2XL U30 ( .A(n2), .B(\u_div/CryTmp[15][1] ), .Y(\u_div/SumTmp[15][1] )
         );
  INVXL U31 ( .A(quotient[14]), .Y(n10) );
  NOR2XL U32 ( .A(\u_div/CryTmp[14][1] ), .B(n10), .Y(n11) );
  NOR2XL U33 ( .A(quotient[14]), .B(n33), .Y(n12) );
  XNOR2XL U34 ( .A(n3), .B(\u_div/CryTmp[13][1] ), .Y(\u_div/SumTmp[13][1] )
         );
  OAI2BB1X2 U35 ( .A0N(n73), .A1N(\u_div/PartRem[15][3] ), .B0(n26), .Y(
        quotient[14]) );
  MXI2X2 U36 ( .A(n43), .B(\u_div/CryTmp[8][1] ), .S0(quotient[8]), .Y(
        \u_div/PartRem[8][1] ) );
  OAI2BB1X2 U37 ( .A0N(n61), .A1N(\u_div/PartRem[9][3] ), .B0(n17), .Y(
        quotient[8]) );
  OAI2BB1X2 U38 ( .A0N(n63), .A1N(\u_div/PartRem[10][3] ), .B0(n16), .Y(
        quotient[9]) );
  MXI2X2 U39 ( .A(n30), .B(\u_div/CryTmp[11][1] ), .S0(quotient[11]), .Y(
        \u_div/PartRem[11][1] ) );
  OAI2BB1X2 U40 ( .A0N(n67), .A1N(\u_div/PartRem[12][3] ), .B0(n14), .Y(
        quotient[11]) );
  OAI2BB1X2 U41 ( .A0N(n69), .A1N(\u_div/PartRem[13][3] ), .B0(n13), .Y(
        quotient[12]) );
  MXI2X2 U42 ( .A(n38), .B(\u_div/CryTmp[3][1] ), .S0(quotient[3]), .Y(
        \u_div/PartRem[3][1] ) );
  OAI2BB1X2 U43 ( .A0N(n51), .A1N(\u_div/PartRem[4][3] ), .B0(n22), .Y(
        quotient[3]) );
  OAI2BB1X2 U44 ( .A0N(n53), .A1N(\u_div/PartRem[5][3] ), .B0(n21), .Y(
        quotient[4]) );
  MXI2XL U45 ( .A(\u_div/PartRem[14][3] ), .B(\u_div/SumTmp[13][3] ), .S0(
        quotient[13]), .Y(n13) );
  MXI2XL U46 ( .A(\u_div/PartRem[13][3] ), .B(\u_div/SumTmp[12][3] ), .S0(
        quotient[12]), .Y(n14) );
  MXI2XL U47 ( .A(\u_div/PartRem[12][3] ), .B(\u_div/SumTmp[11][3] ), .S0(
        quotient[11]), .Y(n15) );
  MXI2XL U48 ( .A(\u_div/PartRem[11][3] ), .B(\u_div/SumTmp[10][3] ), .S0(
        quotient[10]), .Y(n16) );
  MXI2XL U49 ( .A(\u_div/PartRem[10][3] ), .B(\u_div/SumTmp[9][3] ), .S0(
        quotient[9]), .Y(n17) );
  MXI2XL U50 ( .A(\u_div/PartRem[9][3] ), .B(\u_div/SumTmp[8][3] ), .S0(
        quotient[8]), .Y(n18) );
  MXI2XL U51 ( .A(\u_div/PartRem[8][3] ), .B(\u_div/SumTmp[7][3] ), .S0(
        quotient[7]), .Y(n19) );
  MXI2XL U52 ( .A(\u_div/PartRem[7][3] ), .B(\u_div/SumTmp[6][3] ), .S0(
        quotient[6]), .Y(n20) );
  MXI2XL U53 ( .A(\u_div/PartRem[6][3] ), .B(\u_div/SumTmp[5][3] ), .S0(
        quotient[5]), .Y(n21) );
  MXI2XL U54 ( .A(\u_div/PartRem[5][3] ), .B(\u_div/SumTmp[4][3] ), .S0(
        quotient[4]), .Y(n22) );
  MXI2XL U55 ( .A(\u_div/PartRem[4][3] ), .B(\u_div/SumTmp[3][3] ), .S0(
        quotient[3]), .Y(n23) );
  MXI2XL U56 ( .A(\u_div/PartRem[3][3] ), .B(\u_div/SumTmp[2][3] ), .S0(
        quotient[2]), .Y(n24) );
  MXI2XL U57 ( .A(\u_div/PartRem[15][3] ), .B(\u_div/SumTmp[14][3] ), .S0(
        quotient[14]), .Y(n25) );
  MXI2XL U58 ( .A(\u_div/PartRem[16][3] ), .B(\u_div/SumTmp[15][3] ), .S0(
        quotient[15]), .Y(n26) );
  INVXL U59 ( .A(\u_div/CryTmp[16][1] ), .Y(n35) );
  MXI2XL U60 ( .A(a[19]), .B(\u_div/SumTmp[16][3] ), .S0(quotient[16]), .Y(n27) );
  INVXL U61 ( .A(\u_div/CryTmp[1][1] ), .Y(n36) );
  MXI2XL U62 ( .A(n36), .B(\u_div/CryTmp[1][1] ), .S0(quotient[1]), .Y(
        \u_div/PartRem[1][1] ) );
  MXI2XL U63 ( .A(\u_div/PartRem[2][3] ), .B(\u_div/SumTmp[1][3] ), .S0(
        quotient[1]), .Y(n28) );
  NAND2X1 U64 ( .A(n28), .B(n45), .Y(quotient[0]) );
  CLKINVX1 U65 ( .A(\u_div/CryTmp[14][1] ), .Y(n33) );
  CLKINVX1 U66 ( .A(\u_div/CryTmp[5][1] ), .Y(n40) );
  CLKINVX1 U67 ( .A(\u_div/CryTmp[4][1] ), .Y(n39) );
  CLKINVX1 U68 ( .A(\u_div/CryTmp[3][1] ), .Y(n38) );
  CLKINVX1 U69 ( .A(\u_div/CryTmp[12][1] ), .Y(n31) );
  CLKINVX1 U70 ( .A(\u_div/CryTmp[6][1] ), .Y(n41) );
  CLKINVX1 U71 ( .A(\u_div/CryTmp[13][1] ), .Y(n32) );
  CLKINVX1 U72 ( .A(\u_div/CryTmp[11][1] ), .Y(n30) );
  CLKINVX1 U73 ( .A(\u_div/CryTmp[10][1] ), .Y(n29) );
  CLKINVX1 U74 ( .A(\u_div/CryTmp[9][1] ), .Y(n44) );
  CLKINVX1 U75 ( .A(\u_div/CryTmp[8][1] ), .Y(n43) );
  CLKINVX1 U76 ( .A(\u_div/CryTmp[7][1] ), .Y(n42) );
  CLKINVX1 U77 ( .A(\u_div/CryTmp[2][1] ), .Y(n37) );
  CLKINVX1 U78 ( .A(\u_div/CryTmp[15][1] ), .Y(n34) );
  OAI211X1 U79 ( .A0(\u_div/PartRem[1][1] ), .A1(\u_div/CryTmp[0][1] ), .B0(
        \u_div/PartRem[1][2] ), .C0(\u_div/PartRem[1][3] ), .Y(n45) );
  NOR2X1 U80 ( .A(\u_div/CryTmp[1][1] ), .B(\u_div/PartRem[2][1] ), .Y(n46) );
  NOR2BX1 U81 ( .AN(\u_div/PartRem[2][2] ), .B(n46), .Y(n47) );
  XNOR2X1 U82 ( .A(\u_div/PartRem[2][1] ), .B(\u_div/CryTmp[1][1] ), .Y(
        \u_div/SumTmp[1][1] ) );
  XNOR2X1 U83 ( .A(\u_div/PartRem[2][2] ), .B(n46), .Y(\u_div/SumTmp[1][2] )
         );
  XOR2X1 U84 ( .A(\u_div/PartRem[2][3] ), .B(n47), .Y(\u_div/SumTmp[1][3] ) );
  NOR2X1 U85 ( .A(\u_div/CryTmp[2][1] ), .B(\u_div/PartRem[3][1] ), .Y(n48) );
  NOR2BX1 U86 ( .AN(\u_div/PartRem[3][2] ), .B(n48), .Y(n49) );
  XNOR2X1 U87 ( .A(\u_div/PartRem[3][1] ), .B(\u_div/CryTmp[2][1] ), .Y(
        \u_div/SumTmp[2][1] ) );
  XNOR2X1 U88 ( .A(\u_div/PartRem[3][2] ), .B(n48), .Y(\u_div/SumTmp[2][2] )
         );
  XOR2X1 U89 ( .A(\u_div/PartRem[3][3] ), .B(n49), .Y(\u_div/SumTmp[2][3] ) );
  NOR2X1 U90 ( .A(\u_div/CryTmp[3][1] ), .B(\u_div/PartRem[4][1] ), .Y(n50) );
  NOR2BX1 U91 ( .AN(\u_div/PartRem[4][2] ), .B(n50), .Y(n51) );
  XNOR2X1 U92 ( .A(\u_div/PartRem[4][1] ), .B(\u_div/CryTmp[3][1] ), .Y(
        \u_div/SumTmp[3][1] ) );
  XNOR2X1 U93 ( .A(\u_div/PartRem[4][2] ), .B(n50), .Y(\u_div/SumTmp[3][2] )
         );
  XOR2X1 U94 ( .A(\u_div/PartRem[4][3] ), .B(n51), .Y(\u_div/SumTmp[3][3] ) );
  NOR2X1 U95 ( .A(\u_div/CryTmp[4][1] ), .B(\u_div/PartRem[5][1] ), .Y(n52) );
  NOR2BX1 U96 ( .AN(\u_div/PartRem[5][2] ), .B(n52), .Y(n53) );
  XNOR2X1 U97 ( .A(\u_div/PartRem[5][1] ), .B(\u_div/CryTmp[4][1] ), .Y(
        \u_div/SumTmp[4][1] ) );
  XNOR2X1 U98 ( .A(\u_div/PartRem[5][2] ), .B(n52), .Y(\u_div/SumTmp[4][2] )
         );
  XOR2X1 U99 ( .A(\u_div/PartRem[5][3] ), .B(n53), .Y(\u_div/SumTmp[4][3] ) );
  NOR2X1 U100 ( .A(\u_div/CryTmp[5][1] ), .B(\u_div/PartRem[6][1] ), .Y(n54)
         );
  NOR2BX1 U101 ( .AN(\u_div/PartRem[6][2] ), .B(n54), .Y(n55) );
  XNOR2X1 U102 ( .A(\u_div/PartRem[6][1] ), .B(\u_div/CryTmp[5][1] ), .Y(
        \u_div/SumTmp[5][1] ) );
  XNOR2X1 U103 ( .A(\u_div/PartRem[6][2] ), .B(n54), .Y(\u_div/SumTmp[5][2] )
         );
  XOR2X1 U104 ( .A(\u_div/PartRem[6][3] ), .B(n55), .Y(\u_div/SumTmp[5][3] )
         );
  NOR2X1 U105 ( .A(\u_div/CryTmp[6][1] ), .B(\u_div/PartRem[7][1] ), .Y(n56)
         );
  NOR2BX1 U106 ( .AN(\u_div/PartRem[7][2] ), .B(n56), .Y(n57) );
  XNOR2X1 U107 ( .A(\u_div/PartRem[7][1] ), .B(\u_div/CryTmp[6][1] ), .Y(
        \u_div/SumTmp[6][1] ) );
  XNOR2X1 U108 ( .A(\u_div/PartRem[7][2] ), .B(n56), .Y(\u_div/SumTmp[6][2] )
         );
  XOR2X1 U109 ( .A(\u_div/PartRem[7][3] ), .B(n57), .Y(\u_div/SumTmp[6][3] )
         );
  NOR2X1 U110 ( .A(\u_div/CryTmp[7][1] ), .B(\u_div/PartRem[8][1] ), .Y(n58)
         );
  NOR2BX1 U111 ( .AN(\u_div/PartRem[8][2] ), .B(n58), .Y(n59) );
  XNOR2X1 U112 ( .A(\u_div/PartRem[8][1] ), .B(\u_div/CryTmp[7][1] ), .Y(
        \u_div/SumTmp[7][1] ) );
  XNOR2X1 U113 ( .A(\u_div/PartRem[8][2] ), .B(n58), .Y(\u_div/SumTmp[7][2] )
         );
  XOR2X1 U114 ( .A(\u_div/PartRem[8][3] ), .B(n59), .Y(\u_div/SumTmp[7][3] )
         );
  NOR2X1 U115 ( .A(\u_div/CryTmp[8][1] ), .B(\u_div/PartRem[9][1] ), .Y(n60)
         );
  NOR2BX1 U116 ( .AN(\u_div/PartRem[9][2] ), .B(n60), .Y(n61) );
  XNOR2X1 U117 ( .A(\u_div/PartRem[9][1] ), .B(\u_div/CryTmp[8][1] ), .Y(
        \u_div/SumTmp[8][1] ) );
  XNOR2X1 U118 ( .A(\u_div/PartRem[9][2] ), .B(n60), .Y(\u_div/SumTmp[8][2] )
         );
  XOR2X1 U119 ( .A(\u_div/PartRem[9][3] ), .B(n61), .Y(\u_div/SumTmp[8][3] )
         );
  NOR2X1 U120 ( .A(\u_div/CryTmp[9][1] ), .B(\u_div/PartRem[10][1] ), .Y(n62)
         );
  NOR2BX1 U121 ( .AN(\u_div/PartRem[10][2] ), .B(n62), .Y(n63) );
  XNOR2X1 U122 ( .A(\u_div/PartRem[10][1] ), .B(\u_div/CryTmp[9][1] ), .Y(
        \u_div/SumTmp[9][1] ) );
  XNOR2X1 U123 ( .A(\u_div/PartRem[10][2] ), .B(n62), .Y(\u_div/SumTmp[9][2] )
         );
  XOR2X1 U124 ( .A(\u_div/PartRem[10][3] ), .B(n63), .Y(\u_div/SumTmp[9][3] )
         );
  NOR2X1 U125 ( .A(\u_div/CryTmp[10][1] ), .B(\u_div/PartRem[11][1] ), .Y(n64)
         );
  NOR2BX1 U126 ( .AN(\u_div/PartRem[11][2] ), .B(n64), .Y(n65) );
  XNOR2X1 U127 ( .A(\u_div/PartRem[11][1] ), .B(\u_div/CryTmp[10][1] ), .Y(
        \u_div/SumTmp[10][1] ) );
  XNOR2X1 U128 ( .A(\u_div/PartRem[11][2] ), .B(n64), .Y(\u_div/SumTmp[10][2] ) );
  XOR2X1 U129 ( .A(\u_div/PartRem[11][3] ), .B(n65), .Y(\u_div/SumTmp[10][3] )
         );
  NOR2X1 U130 ( .A(\u_div/CryTmp[11][1] ), .B(\u_div/PartRem[12][1] ), .Y(n66)
         );
  NOR2BX1 U131 ( .AN(\u_div/PartRem[12][2] ), .B(n66), .Y(n67) );
  XNOR2X1 U132 ( .A(\u_div/PartRem[12][1] ), .B(\u_div/CryTmp[11][1] ), .Y(
        \u_div/SumTmp[11][1] ) );
  XNOR2X1 U133 ( .A(\u_div/PartRem[12][2] ), .B(n66), .Y(\u_div/SumTmp[11][2] ) );
  XOR2X1 U134 ( .A(\u_div/PartRem[12][3] ), .B(n67), .Y(\u_div/SumTmp[11][3] )
         );
  NOR2X1 U135 ( .A(\u_div/CryTmp[12][1] ), .B(n1), .Y(n68) );
  NOR2BX1 U136 ( .AN(\u_div/PartRem[13][2] ), .B(n68), .Y(n69) );
  XNOR2X1 U137 ( .A(\u_div/PartRem[13][2] ), .B(n68), .Y(\u_div/SumTmp[12][2] ) );
  XOR2X1 U138 ( .A(\u_div/PartRem[13][3] ), .B(n69), .Y(\u_div/SumTmp[12][3] )
         );
  NOR2X1 U139 ( .A(\u_div/CryTmp[13][1] ), .B(n3), .Y(n70) );
  NOR2BX1 U140 ( .AN(\u_div/PartRem[14][2] ), .B(n70), .Y(n71) );
  XNOR2X1 U141 ( .A(\u_div/PartRem[14][2] ), .B(n70), .Y(\u_div/SumTmp[13][2] ) );
  XOR2X1 U142 ( .A(\u_div/PartRem[14][3] ), .B(n71), .Y(\u_div/SumTmp[13][3] )
         );
  NOR2X1 U143 ( .A(\u_div/CryTmp[14][1] ), .B(\u_div/PartRem[15][1] ), .Y(n72)
         );
  NOR2BX1 U144 ( .AN(\u_div/PartRem[15][2] ), .B(n72), .Y(n73) );
  XNOR2X1 U145 ( .A(\u_div/PartRem[15][1] ), .B(\u_div/CryTmp[14][1] ), .Y(
        \u_div/SumTmp[14][1] ) );
  XNOR2X1 U146 ( .A(\u_div/PartRem[15][2] ), .B(n72), .Y(\u_div/SumTmp[14][2] ) );
  XOR2X1 U147 ( .A(\u_div/PartRem[15][3] ), .B(n73), .Y(\u_div/SumTmp[14][3] )
         );
  NOR2X1 U148 ( .A(\u_div/CryTmp[15][1] ), .B(n2), .Y(n74) );
  NOR2BX1 U149 ( .AN(\u_div/PartRem[16][2] ), .B(n74), .Y(n75) );
  XNOR2X1 U150 ( .A(\u_div/PartRem[16][2] ), .B(n74), .Y(\u_div/SumTmp[15][2] ) );
  NOR2X1 U151 ( .A(\u_div/CryTmp[16][1] ), .B(\u_div/CryTmp[17][1] ), .Y(n76)
         );
  NOR2BX1 U152 ( .AN(\u_div/CryTmp[18][1] ), .B(n76), .Y(n77) );
  XNOR2X1 U153 ( .A(\u_div/CryTmp[17][1] ), .B(\u_div/CryTmp[16][1] ), .Y(
        \u_div/SumTmp[16][1] ) );
  XNOR2X1 U154 ( .A(\u_div/CryTmp[18][1] ), .B(n76), .Y(\u_div/SumTmp[16][2] )
         );
  XOR2X1 U155 ( .A(a[19]), .B(n77), .Y(\u_div/SumTmp[16][3] ) );
endmodule


module CONT_DW_div_uns_9 ( a, b, quotient, remainder, divide_by_0 );
  input [19:0] a;
  input [8:0] b;
  output [19:0] quotient;
  output [8:0] remainder;
  output divide_by_0;
  wire   n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         \u_div/SumTmp[1][2] , \u_div/SumTmp[1][3] , \u_div/SumTmp[1][4] ,
         \u_div/SumTmp[1][5] , \u_div/SumTmp[1][6] , \u_div/SumTmp[1][7] ,
         \u_div/SumTmp[1][8] , \u_div/SumTmp[2][1] , \u_div/SumTmp[2][2] ,
         \u_div/SumTmp[2][3] , \u_div/SumTmp[2][4] , \u_div/SumTmp[2][5] ,
         \u_div/SumTmp[2][6] , \u_div/SumTmp[2][7] , \u_div/SumTmp[2][8] ,
         \u_div/SumTmp[3][0] , \u_div/SumTmp[3][1] , \u_div/SumTmp[3][2] ,
         \u_div/SumTmp[3][3] , \u_div/SumTmp[3][4] , \u_div/SumTmp[3][5] ,
         \u_div/SumTmp[3][6] , \u_div/SumTmp[3][7] , \u_div/SumTmp[3][8] ,
         \u_div/SumTmp[4][0] , \u_div/SumTmp[4][1] , \u_div/SumTmp[4][2] ,
         \u_div/SumTmp[4][3] , \u_div/SumTmp[4][4] , \u_div/SumTmp[4][5] ,
         \u_div/SumTmp[4][6] , \u_div/SumTmp[4][7] , \u_div/SumTmp[4][8] ,
         \u_div/SumTmp[5][0] , \u_div/SumTmp[5][1] , \u_div/SumTmp[5][2] ,
         \u_div/SumTmp[5][3] , \u_div/SumTmp[5][4] , \u_div/SumTmp[5][5] ,
         \u_div/SumTmp[5][6] , \u_div/SumTmp[5][7] , \u_div/SumTmp[5][8] ,
         \u_div/SumTmp[6][0] , \u_div/SumTmp[6][1] , \u_div/SumTmp[6][2] ,
         \u_div/SumTmp[6][3] , \u_div/SumTmp[6][4] , \u_div/SumTmp[6][5] ,
         \u_div/SumTmp[6][6] , \u_div/SumTmp[6][7] , \u_div/SumTmp[6][8] ,
         \u_div/SumTmp[7][0] , \u_div/SumTmp[7][1] , \u_div/SumTmp[7][2] ,
         \u_div/SumTmp[7][3] , \u_div/SumTmp[7][4] , \u_div/SumTmp[7][5] ,
         \u_div/SumTmp[7][6] , \u_div/SumTmp[7][7] , \u_div/SumTmp[7][8] ,
         \u_div/SumTmp[8][0] , \u_div/SumTmp[8][1] , \u_div/SumTmp[8][2] ,
         \u_div/SumTmp[8][3] , \u_div/SumTmp[8][4] , \u_div/SumTmp[8][5] ,
         \u_div/SumTmp[8][6] , \u_div/SumTmp[8][7] , \u_div/SumTmp[8][8] ,
         \u_div/SumTmp[9][0] , \u_div/SumTmp[9][1] , \u_div/SumTmp[9][2] ,
         \u_div/SumTmp[9][3] , \u_div/SumTmp[9][4] , \u_div/SumTmp[9][5] ,
         \u_div/SumTmp[9][6] , \u_div/SumTmp[9][7] , \u_div/SumTmp[9][8] ,
         \u_div/SumTmp[10][0] , \u_div/SumTmp[10][1] , \u_div/SumTmp[10][2] ,
         \u_div/SumTmp[10][3] , \u_div/SumTmp[10][4] , \u_div/SumTmp[10][5] ,
         \u_div/SumTmp[10][6] , \u_div/SumTmp[10][7] , \u_div/SumTmp[10][8] ,
         \u_div/SumTmp[11][0] , \u_div/SumTmp[11][1] , \u_div/SumTmp[11][2] ,
         \u_div/SumTmp[11][3] , \u_div/SumTmp[11][4] , \u_div/SumTmp[11][5] ,
         \u_div/SumTmp[11][6] , \u_div/SumTmp[11][7] , \u_div/SumTmp[11][8] ,
         \u_div/SumTmp[14][0] , \u_div/SumTmp[15][0] , \u_div/SumTmp[16][0] ,
         \u_div/SumTmp[17][0] , \u_div/SumTmp[18][0] , \u_div/SumTmp[19][0] ,
         \u_div/PartRem[1][6] , \u_div/PartRem[1][7] , \u_div/PartRem[1][8] ,
         \u_div/PartRem[1][9] , \u_div/PartRem[2][3] , \u_div/PartRem[2][4] ,
         \u_div/PartRem[2][5] , \u_div/PartRem[2][6] , \u_div/PartRem[2][7] ,
         \u_div/PartRem[2][8] , \u_div/PartRem[2][9] , \u_div/PartRem[3][3] ,
         \u_div/PartRem[3][4] , \u_div/PartRem[3][5] , \u_div/PartRem[3][6] ,
         \u_div/PartRem[3][7] , \u_div/PartRem[3][8] , \u_div/PartRem[3][9] ,
         \u_div/PartRem[4][3] , \u_div/PartRem[4][4] , \u_div/PartRem[4][5] ,
         \u_div/PartRem[4][6] , \u_div/PartRem[4][7] , \u_div/PartRem[4][8] ,
         \u_div/PartRem[4][9] , \u_div/PartRem[5][3] , \u_div/PartRem[5][4] ,
         \u_div/PartRem[5][5] , \u_div/PartRem[5][6] , \u_div/PartRem[5][7] ,
         \u_div/PartRem[5][8] , \u_div/PartRem[5][9] , \u_div/PartRem[6][3] ,
         \u_div/PartRem[6][4] , \u_div/PartRem[6][5] , \u_div/PartRem[6][6] ,
         \u_div/PartRem[6][7] , \u_div/PartRem[6][8] , \u_div/PartRem[6][9] ,
         \u_div/PartRem[7][3] , \u_div/PartRem[7][4] , \u_div/PartRem[7][5] ,
         \u_div/PartRem[7][6] , \u_div/PartRem[7][7] , \u_div/PartRem[7][8] ,
         \u_div/PartRem[7][9] , \u_div/PartRem[8][3] , \u_div/PartRem[8][4] ,
         \u_div/PartRem[8][5] , \u_div/PartRem[8][6] , \u_div/PartRem[8][7] ,
         \u_div/PartRem[8][8] , \u_div/PartRem[8][9] , \u_div/PartRem[9][3] ,
         \u_div/PartRem[9][4] , \u_div/PartRem[9][5] , \u_div/PartRem[9][6] ,
         \u_div/PartRem[9][7] , \u_div/PartRem[9][8] , \u_div/PartRem[9][9] ,
         \u_div/PartRem[10][3] , \u_div/PartRem[10][4] ,
         \u_div/PartRem[10][5] , \u_div/PartRem[10][6] ,
         \u_div/PartRem[10][7] , \u_div/PartRem[10][8] ,
         \u_div/PartRem[10][9] , \u_div/PartRem[11][3] ,
         \u_div/PartRem[11][4] , \u_div/PartRem[11][5] ,
         \u_div/PartRem[11][6] , \u_div/PartRem[11][7] ,
         \u_div/PartRem[11][8] , \u_div/PartRem[11][9] ,
         \u_div/u_add_PartRem_0_1/n6 , \u_div/u_add_PartRem_0_1/n5 ,
         \u_div/u_add_PartRem_0_1/n3 , \u_div/u_add_PartRem_0_1/n2 ,
         \u_div/u_add_PartRem_0_2/n6 , \u_div/u_add_PartRem_0_2/n5 ,
         \u_div/u_add_PartRem_0_2/n3 , \u_div/u_add_PartRem_0_2/n2 ,
         \u_div/u_add_PartRem_0_3/n6 , \u_div/u_add_PartRem_0_3/n5 ,
         \u_div/u_add_PartRem_0_3/n3 , \u_div/u_add_PartRem_0_3/n2 ,
         \u_div/u_add_PartRem_0_4/n6 , \u_div/u_add_PartRem_0_4/n5 ,
         \u_div/u_add_PartRem_0_4/n3 , \u_div/u_add_PartRem_0_4/n2 ,
         \u_div/u_add_PartRem_0_5/n6 , \u_div/u_add_PartRem_0_5/n5 ,
         \u_div/u_add_PartRem_0_5/n3 , \u_div/u_add_PartRem_0_5/n2 ,
         \u_div/u_add_PartRem_0_6/n6 , \u_div/u_add_PartRem_0_6/n5 ,
         \u_div/u_add_PartRem_0_6/n3 , \u_div/u_add_PartRem_0_6/n2 ,
         \u_div/u_add_PartRem_0_7/n6 , \u_div/u_add_PartRem_0_7/n5 ,
         \u_div/u_add_PartRem_0_7/n3 , \u_div/u_add_PartRem_0_7/n2 ,
         \u_div/u_add_PartRem_0_8/n6 , \u_div/u_add_PartRem_0_8/n5 ,
         \u_div/u_add_PartRem_0_8/n3 , \u_div/u_add_PartRem_0_8/n2 ,
         \u_div/u_add_PartRem_0_9/n6 , \u_div/u_add_PartRem_0_9/n5 ,
         \u_div/u_add_PartRem_0_9/n3 , \u_div/u_add_PartRem_0_9/n2 ,
         \u_div/u_add_PartRem_0_10/n6 , \u_div/u_add_PartRem_0_10/n5 ,
         \u_div/u_add_PartRem_0_10/n3 , \u_div/u_add_PartRem_0_10/n2 ,
         \u_div/u_add_PartRem_1_11/n5 , \u_div/u_add_PartRem_1_11/n4 ,
         \u_div/u_add_PartRem_1_11/n2 , n1, n2, n3, n4, n5, n6, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign \u_div/SumTmp[3][0]  = a[3];
  assign \u_div/SumTmp[4][0]  = a[4];
  assign \u_div/SumTmp[5][0]  = a[5];
  assign \u_div/SumTmp[6][0]  = a[6];
  assign \u_div/SumTmp[7][0]  = a[7];
  assign \u_div/SumTmp[8][0]  = a[8];
  assign \u_div/SumTmp[9][0]  = a[9];
  assign \u_div/SumTmp[10][0]  = a[10];
  assign \u_div/SumTmp[11][0]  = a[11];
  assign \u_div/SumTmp[11][1]  = a[12];
  assign \u_div/SumTmp[11][2]  = a[13];
  assign \u_div/SumTmp[14][0]  = a[14];
  assign \u_div/SumTmp[15][0]  = a[15];
  assign \u_div/SumTmp[16][0]  = a[16];
  assign \u_div/SumTmp[17][0]  = a[17];
  assign \u_div/SumTmp[18][0]  = a[18];
  assign \u_div/SumTmp[19][0]  = a[19];

  ADDHXL \u_div/u_add_PartRem_0_1/U9  ( .A(\u_div/PartRem[2][4] ), .B(
        \u_div/PartRem[2][3] ), .CO(\u_div/u_add_PartRem_0_1/n6 ), .S(
        \u_div/SumTmp[1][4] ) );
  ADDHXL \u_div/u_add_PartRem_0_1/U8  ( .A(\u_div/PartRem[2][5] ), .B(
        \u_div/u_add_PartRem_0_1/n6 ), .CO(\u_div/u_add_PartRem_0_1/n5 ), .S(
        \u_div/SumTmp[1][5] ) );
  ADDHXL \u_div/u_add_PartRem_0_1/U3  ( .A(\u_div/PartRem[2][8] ), .B(
        \u_div/u_add_PartRem_0_1/n3 ), .CO(\u_div/u_add_PartRem_0_1/n2 ), .S(
        \u_div/SumTmp[1][8] ) );
  ADDHXL \u_div/u_add_PartRem_0_2/U9  ( .A(\u_div/PartRem[3][4] ), .B(
        \u_div/PartRem[3][3] ), .CO(\u_div/u_add_PartRem_0_2/n6 ), .S(
        \u_div/SumTmp[2][4] ) );
  ADDHXL \u_div/u_add_PartRem_0_2/U8  ( .A(\u_div/PartRem[3][5] ), .B(
        \u_div/u_add_PartRem_0_2/n6 ), .CO(\u_div/u_add_PartRem_0_2/n5 ), .S(
        \u_div/SumTmp[2][5] ) );
  ADDHXL \u_div/u_add_PartRem_0_2/U3  ( .A(\u_div/PartRem[3][8] ), .B(
        \u_div/u_add_PartRem_0_2/n3 ), .CO(\u_div/u_add_PartRem_0_2/n2 ), .S(
        \u_div/SumTmp[2][8] ) );
  ADDHXL \u_div/u_add_PartRem_0_3/U9  ( .A(\u_div/PartRem[4][4] ), .B(
        \u_div/PartRem[4][3] ), .CO(\u_div/u_add_PartRem_0_3/n6 ), .S(
        \u_div/SumTmp[3][4] ) );
  ADDHXL \u_div/u_add_PartRem_0_3/U8  ( .A(\u_div/PartRem[4][5] ), .B(
        \u_div/u_add_PartRem_0_3/n6 ), .CO(\u_div/u_add_PartRem_0_3/n5 ), .S(
        \u_div/SumTmp[3][5] ) );
  ADDHXL \u_div/u_add_PartRem_0_3/U3  ( .A(\u_div/PartRem[4][8] ), .B(
        \u_div/u_add_PartRem_0_3/n3 ), .CO(\u_div/u_add_PartRem_0_3/n2 ), .S(
        \u_div/SumTmp[3][8] ) );
  ADDHXL \u_div/u_add_PartRem_0_4/U9  ( .A(\u_div/PartRem[5][4] ), .B(
        \u_div/PartRem[5][3] ), .CO(\u_div/u_add_PartRem_0_4/n6 ), .S(
        \u_div/SumTmp[4][4] ) );
  ADDHXL \u_div/u_add_PartRem_0_4/U8  ( .A(\u_div/PartRem[5][5] ), .B(
        \u_div/u_add_PartRem_0_4/n6 ), .CO(\u_div/u_add_PartRem_0_4/n5 ), .S(
        \u_div/SumTmp[4][5] ) );
  ADDHXL \u_div/u_add_PartRem_0_4/U3  ( .A(\u_div/PartRem[5][8] ), .B(
        \u_div/u_add_PartRem_0_4/n3 ), .CO(\u_div/u_add_PartRem_0_4/n2 ), .S(
        \u_div/SumTmp[4][8] ) );
  ADDHXL \u_div/u_add_PartRem_0_5/U9  ( .A(\u_div/PartRem[6][4] ), .B(
        \u_div/PartRem[6][3] ), .CO(\u_div/u_add_PartRem_0_5/n6 ), .S(
        \u_div/SumTmp[5][4] ) );
  ADDHXL \u_div/u_add_PartRem_0_5/U8  ( .A(\u_div/PartRem[6][5] ), .B(
        \u_div/u_add_PartRem_0_5/n6 ), .CO(\u_div/u_add_PartRem_0_5/n5 ), .S(
        \u_div/SumTmp[5][5] ) );
  ADDHXL \u_div/u_add_PartRem_0_5/U3  ( .A(\u_div/PartRem[6][8] ), .B(
        \u_div/u_add_PartRem_0_5/n3 ), .CO(\u_div/u_add_PartRem_0_5/n2 ), .S(
        \u_div/SumTmp[5][8] ) );
  ADDHXL \u_div/u_add_PartRem_0_6/U9  ( .A(\u_div/PartRem[7][4] ), .B(
        \u_div/PartRem[7][3] ), .CO(\u_div/u_add_PartRem_0_6/n6 ), .S(
        \u_div/SumTmp[6][4] ) );
  ADDHXL \u_div/u_add_PartRem_0_6/U8  ( .A(\u_div/PartRem[7][5] ), .B(
        \u_div/u_add_PartRem_0_6/n6 ), .CO(\u_div/u_add_PartRem_0_6/n5 ), .S(
        \u_div/SumTmp[6][5] ) );
  ADDHXL \u_div/u_add_PartRem_0_6/U3  ( .A(\u_div/PartRem[7][8] ), .B(
        \u_div/u_add_PartRem_0_6/n3 ), .CO(\u_div/u_add_PartRem_0_6/n2 ), .S(
        \u_div/SumTmp[6][8] ) );
  ADDHXL \u_div/u_add_PartRem_0_7/U9  ( .A(\u_div/PartRem[8][4] ), .B(
        \u_div/PartRem[8][3] ), .CO(\u_div/u_add_PartRem_0_7/n6 ), .S(
        \u_div/SumTmp[7][4] ) );
  ADDHXL \u_div/u_add_PartRem_0_7/U8  ( .A(\u_div/PartRem[8][5] ), .B(
        \u_div/u_add_PartRem_0_7/n6 ), .CO(\u_div/u_add_PartRem_0_7/n5 ), .S(
        \u_div/SumTmp[7][5] ) );
  ADDHXL \u_div/u_add_PartRem_0_7/U3  ( .A(\u_div/PartRem[8][8] ), .B(
        \u_div/u_add_PartRem_0_7/n3 ), .CO(\u_div/u_add_PartRem_0_7/n2 ), .S(
        \u_div/SumTmp[7][8] ) );
  ADDHXL \u_div/u_add_PartRem_0_8/U9  ( .A(\u_div/PartRem[9][4] ), .B(
        \u_div/PartRem[9][3] ), .CO(\u_div/u_add_PartRem_0_8/n6 ), .S(
        \u_div/SumTmp[8][4] ) );
  ADDHXL \u_div/u_add_PartRem_0_8/U8  ( .A(\u_div/PartRem[9][5] ), .B(
        \u_div/u_add_PartRem_0_8/n6 ), .CO(\u_div/u_add_PartRem_0_8/n5 ), .S(
        \u_div/SumTmp[8][5] ) );
  ADDHXL \u_div/u_add_PartRem_0_8/U3  ( .A(\u_div/PartRem[9][8] ), .B(
        \u_div/u_add_PartRem_0_8/n3 ), .CO(\u_div/u_add_PartRem_0_8/n2 ), .S(
        \u_div/SumTmp[8][8] ) );
  ADDHXL \u_div/u_add_PartRem_0_9/U9  ( .A(\u_div/PartRem[10][4] ), .B(
        \u_div/PartRem[10][3] ), .CO(\u_div/u_add_PartRem_0_9/n6 ), .S(
        \u_div/SumTmp[9][4] ) );
  ADDHXL \u_div/u_add_PartRem_0_9/U8  ( .A(\u_div/PartRem[10][5] ), .B(
        \u_div/u_add_PartRem_0_9/n6 ), .CO(\u_div/u_add_PartRem_0_9/n5 ), .S(
        \u_div/SumTmp[9][5] ) );
  ADDHXL \u_div/u_add_PartRem_0_9/U3  ( .A(\u_div/PartRem[10][8] ), .B(
        \u_div/u_add_PartRem_0_9/n3 ), .CO(\u_div/u_add_PartRem_0_9/n2 ), .S(
        \u_div/SumTmp[9][8] ) );
  ADDHXL \u_div/u_add_PartRem_0_10/U9  ( .A(\u_div/PartRem[11][4] ), .B(
        \u_div/PartRem[11][3] ), .CO(\u_div/u_add_PartRem_0_10/n6 ), .S(
        \u_div/SumTmp[10][4] ) );
  ADDHXL \u_div/u_add_PartRem_0_10/U8  ( .A(\u_div/PartRem[11][5] ), .B(
        \u_div/u_add_PartRem_0_10/n6 ), .CO(\u_div/u_add_PartRem_0_10/n5 ), 
        .S(\u_div/SumTmp[10][5] ) );
  ADDHXL \u_div/u_add_PartRem_0_10/U3  ( .A(\u_div/PartRem[11][8] ), .B(
        \u_div/u_add_PartRem_0_10/n3 ), .CO(\u_div/u_add_PartRem_0_10/n2 ), 
        .S(\u_div/SumTmp[10][8] ) );
  ADDHXL \u_div/u_add_PartRem_1_11/U8  ( .A(\u_div/SumTmp[15][0] ), .B(
        \u_div/SumTmp[14][0] ), .CO(\u_div/u_add_PartRem_1_11/n5 ), .S(
        \u_div/SumTmp[11][4] ) );
  ADDHXL \u_div/u_add_PartRem_1_11/U7  ( .A(\u_div/SumTmp[16][0] ), .B(
        \u_div/u_add_PartRem_1_11/n5 ), .CO(\u_div/u_add_PartRem_1_11/n4 ), 
        .S(\u_div/SumTmp[11][5] ) );
  MX2XL \u_div/u_mx_PartRem_0_3_0  ( .A(\u_div/SumTmp[3][0] ), .B(
        \u_div/SumTmp[3][0] ), .S0(quotient[3]), .Y(\u_div/SumTmp[2][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_2_1  ( .A(\u_div/SumTmp[2][1] ), .B(
        \u_div/SumTmp[2][1] ), .S0(quotient[2]), .Y(\u_div/SumTmp[1][2] ) );
  MX2XL \u_div/u_mx_PartRem_0_11_7  ( .A(\u_div/SumTmp[18][0] ), .B(
        \u_div/SumTmp[11][7] ), .S0(n4), .Y(\u_div/PartRem[11][8] ) );
  MX2X1 \u_div/u_mx_PartRem_0_11_6  ( .A(\u_div/SumTmp[17][0] ), .B(
        \u_div/SumTmp[11][6] ), .S0(n4), .Y(\u_div/PartRem[11][7] ) );
  MX2X1 \u_div/u_mx_PartRem_0_11_5  ( .A(\u_div/SumTmp[16][0] ), .B(
        \u_div/SumTmp[11][5] ), .S0(n4), .Y(\u_div/PartRem[11][6] ) );
  MX2XL \u_div/u_mx_PartRem_0_11_8  ( .A(\u_div/SumTmp[19][0] ), .B(
        \u_div/SumTmp[11][8] ), .S0(n4), .Y(\u_div/PartRem[11][9] ) );
  MX2XL \u_div/u_mx_PartRem_0_11_4  ( .A(\u_div/SumTmp[15][0] ), .B(
        \u_div/SumTmp[11][4] ), .S0(n4), .Y(\u_div/PartRem[11][5] ) );
  MX2XL \u_div/u_mx_PartRem_0_5_0  ( .A(\u_div/SumTmp[5][0] ), .B(
        \u_div/SumTmp[5][0] ), .S0(quotient[5]), .Y(\u_div/SumTmp[4][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_4_1  ( .A(\u_div/SumTmp[4][1] ), .B(
        \u_div/SumTmp[4][1] ), .S0(quotient[4]), .Y(\u_div/SumTmp[3][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_3_2  ( .A(\u_div/SumTmp[3][2] ), .B(
        \u_div/SumTmp[3][2] ), .S0(quotient[3]), .Y(\u_div/PartRem[3][3] ) );
  MX2XL \u_div/u_mx_PartRem_0_6_0  ( .A(\u_div/SumTmp[6][0] ), .B(
        \u_div/SumTmp[6][0] ), .S0(quotient[6]), .Y(\u_div/SumTmp[5][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_5_1  ( .A(\u_div/SumTmp[5][1] ), .B(
        \u_div/SumTmp[5][1] ), .S0(quotient[5]), .Y(\u_div/SumTmp[4][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_4_2  ( .A(\u_div/SumTmp[4][2] ), .B(
        \u_div/SumTmp[4][2] ), .S0(quotient[4]), .Y(\u_div/PartRem[4][3] ) );
  MX2XL \u_div/u_mx_PartRem_0_7_0  ( .A(\u_div/SumTmp[7][0] ), .B(
        \u_div/SumTmp[7][0] ), .S0(quotient[7]), .Y(\u_div/SumTmp[6][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_6_1  ( .A(\u_div/SumTmp[6][1] ), .B(
        \u_div/SumTmp[6][1] ), .S0(quotient[6]), .Y(\u_div/SumTmp[5][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_5_2  ( .A(\u_div/SumTmp[5][2] ), .B(
        \u_div/SumTmp[5][2] ), .S0(quotient[5]), .Y(\u_div/PartRem[5][3] ) );
  MX2XL \u_div/u_mx_PartRem_0_8_0  ( .A(\u_div/SumTmp[8][0] ), .B(
        \u_div/SumTmp[8][0] ), .S0(quotient[8]), .Y(\u_div/SumTmp[7][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_7_1  ( .A(\u_div/SumTmp[7][1] ), .B(
        \u_div/SumTmp[7][1] ), .S0(quotient[7]), .Y(\u_div/SumTmp[6][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_6_2  ( .A(\u_div/SumTmp[6][2] ), .B(
        \u_div/SumTmp[6][2] ), .S0(quotient[6]), .Y(\u_div/PartRem[6][3] ) );
  MX2XL \u_div/u_mx_PartRem_0_9_0  ( .A(\u_div/SumTmp[9][0] ), .B(
        \u_div/SumTmp[9][0] ), .S0(n6), .Y(\u_div/SumTmp[8][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_8_1  ( .A(\u_div/SumTmp[8][1] ), .B(
        \u_div/SumTmp[8][1] ), .S0(quotient[8]), .Y(\u_div/SumTmp[7][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_7_2  ( .A(\u_div/SumTmp[7][2] ), .B(
        \u_div/SumTmp[7][2] ), .S0(quotient[7]), .Y(\u_div/PartRem[7][3] ) );
  MX2XL \u_div/u_mx_PartRem_0_10_0  ( .A(\u_div/SumTmp[10][0] ), .B(
        \u_div/SumTmp[10][0] ), .S0(n5), .Y(\u_div/SumTmp[9][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_9_1  ( .A(\u_div/SumTmp[9][1] ), .B(
        \u_div/SumTmp[9][1] ), .S0(n6), .Y(\u_div/SumTmp[8][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_8_2  ( .A(\u_div/SumTmp[8][2] ), .B(
        \u_div/SumTmp[8][2] ), .S0(quotient[8]), .Y(\u_div/PartRem[8][3] ) );
  MX2XL \u_div/u_mx_PartRem_0_4_0  ( .A(\u_div/SumTmp[4][0] ), .B(
        \u_div/SumTmp[4][0] ), .S0(quotient[4]), .Y(\u_div/SumTmp[3][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_3_1  ( .A(\u_div/SumTmp[3][1] ), .B(
        \u_div/SumTmp[3][1] ), .S0(quotient[3]), .Y(\u_div/SumTmp[2][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_2_2  ( .A(\u_div/SumTmp[2][2] ), .B(
        \u_div/SumTmp[2][2] ), .S0(quotient[2]), .Y(\u_div/PartRem[2][3] ) );
  MX2XL \u_div/u_mx_PartRem_0_11_0  ( .A(\u_div/SumTmp[11][0] ), .B(
        \u_div/SumTmp[11][0] ), .S0(n4), .Y(\u_div/SumTmp[10][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_10_1  ( .A(\u_div/SumTmp[10][1] ), .B(
        \u_div/SumTmp[10][1] ), .S0(n5), .Y(\u_div/SumTmp[9][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_9_2  ( .A(\u_div/SumTmp[9][2] ), .B(
        \u_div/SumTmp[9][2] ), .S0(n6), .Y(\u_div/PartRem[9][3] ) );
  MX2XL \u_div/u_mx_PartRem_0_11_1  ( .A(\u_div/SumTmp[11][1] ), .B(
        \u_div/SumTmp[11][1] ), .S0(n4), .Y(\u_div/SumTmp[10][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_10_2  ( .A(\u_div/SumTmp[10][2] ), .B(
        \u_div/SumTmp[10][2] ), .S0(n5), .Y(\u_div/PartRem[10][3] ) );
  MX2X1 \u_div/u_mx_PartRem_0_11_2  ( .A(\u_div/SumTmp[11][2] ), .B(
        \u_div/SumTmp[11][2] ), .S0(n4), .Y(\u_div/PartRem[11][3] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_10_7  ( .A(\u_div/PartRem[11][7] ), .B(
        \u_div/SumTmp[10][7] ), .S0(n5), .Y(\u_div/PartRem[10][8] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_10_6  ( .A(\u_div/PartRem[11][6] ), .B(
        \u_div/SumTmp[10][6] ), .S0(n5), .Y(\u_div/PartRem[10][7] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_10_5  ( .A(\u_div/PartRem[11][5] ), .B(
        \u_div/SumTmp[10][5] ), .S0(n5), .Y(\u_div/PartRem[10][6] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_10_8  ( .A(\u_div/PartRem[11][8] ), .B(
        \u_div/SumTmp[10][8] ), .S0(n5), .Y(\u_div/PartRem[10][9] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_3_3  ( .A(\u_div/PartRem[4][3] ), .B(
        \u_div/SumTmp[3][3] ), .S0(quotient[3]), .Y(\u_div/PartRem[3][4] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_4_3  ( .A(\u_div/PartRem[5][3] ), .B(
        \u_div/SumTmp[4][3] ), .S0(quotient[4]), .Y(\u_div/PartRem[4][4] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_5_3  ( .A(\u_div/PartRem[6][3] ), .B(
        \u_div/SumTmp[5][3] ), .S0(quotient[5]), .Y(\u_div/PartRem[5][4] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_6_3  ( .A(\u_div/PartRem[7][3] ), .B(
        \u_div/SumTmp[6][3] ), .S0(quotient[6]), .Y(\u_div/PartRem[6][4] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_7_3  ( .A(\u_div/PartRem[8][3] ), .B(
        \u_div/SumTmp[7][3] ), .S0(quotient[7]), .Y(\u_div/PartRem[7][4] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_8_3  ( .A(\u_div/PartRem[9][3] ), .B(
        \u_div/SumTmp[8][3] ), .S0(quotient[8]), .Y(\u_div/PartRem[8][4] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_2_3  ( .A(\u_div/PartRem[3][3] ), .B(
        \u_div/SumTmp[2][3] ), .S0(quotient[2]), .Y(\u_div/PartRem[2][4] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_9_3  ( .A(\u_div/PartRem[10][3] ), .B(
        \u_div/SumTmp[9][3] ), .S0(n6), .Y(\u_div/PartRem[9][4] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_10_3  ( .A(\u_div/PartRem[11][3] ), .B(
        \u_div/SumTmp[10][3] ), .S0(n5), .Y(\u_div/PartRem[10][4] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_10_4  ( .A(\u_div/PartRem[11][4] ), .B(
        \u_div/SumTmp[10][4] ), .S0(n5), .Y(\u_div/PartRem[10][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_9_7  ( .A(\u_div/PartRem[10][7] ), .B(
        \u_div/SumTmp[9][7] ), .S0(n6), .Y(\u_div/PartRem[9][8] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_9_6  ( .A(\u_div/PartRem[10][6] ), .B(
        \u_div/SumTmp[9][6] ), .S0(n6), .Y(\u_div/PartRem[9][7] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_9_5  ( .A(\u_div/PartRem[10][5] ), .B(
        \u_div/SumTmp[9][5] ), .S0(n6), .Y(\u_div/PartRem[9][6] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_9_8  ( .A(\u_div/PartRem[10][8] ), .B(
        \u_div/SumTmp[9][8] ), .S0(n6), .Y(\u_div/PartRem[9][9] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_2_4  ( .A(\u_div/PartRem[3][4] ), .B(
        \u_div/SumTmp[2][4] ), .S0(quotient[2]), .Y(\u_div/PartRem[2][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_3_4  ( .A(\u_div/PartRem[4][4] ), .B(
        \u_div/SumTmp[3][4] ), .S0(quotient[3]), .Y(\u_div/PartRem[3][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_4_4  ( .A(\u_div/PartRem[5][4] ), .B(
        \u_div/SumTmp[4][4] ), .S0(quotient[4]), .Y(\u_div/PartRem[4][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_5_4  ( .A(\u_div/PartRem[6][4] ), .B(
        \u_div/SumTmp[5][4] ), .S0(quotient[5]), .Y(\u_div/PartRem[5][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_6_4  ( .A(\u_div/PartRem[7][4] ), .B(
        \u_div/SumTmp[6][4] ), .S0(quotient[6]), .Y(\u_div/PartRem[6][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_7_4  ( .A(\u_div/PartRem[8][4] ), .B(
        \u_div/SumTmp[7][4] ), .S0(quotient[7]), .Y(\u_div/PartRem[7][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_8_4  ( .A(\u_div/PartRem[9][4] ), .B(
        \u_div/SumTmp[8][4] ), .S0(quotient[8]), .Y(\u_div/PartRem[8][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_9_4  ( .A(\u_div/PartRem[10][4] ), .B(
        \u_div/SumTmp[9][4] ), .S0(n6), .Y(\u_div/PartRem[9][5] ) );
  MX2XL \u_div/u_mx_PartRem_0_1_7  ( .A(\u_div/PartRem[2][7] ), .B(
        \u_div/SumTmp[1][7] ), .S0(quotient[1]), .Y(\u_div/PartRem[1][8] ) );
  MX2XL \u_div/u_mx_PartRem_0_1_8  ( .A(\u_div/PartRem[2][8] ), .B(
        \u_div/SumTmp[1][8] ), .S0(quotient[1]), .Y(\u_div/PartRem[1][9] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_8_7  ( .A(\u_div/PartRem[9][7] ), .B(
        \u_div/SumTmp[8][7] ), .S0(quotient[8]), .Y(\u_div/PartRem[8][8] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_2_6  ( .A(\u_div/PartRem[3][6] ), .B(
        \u_div/SumTmp[2][6] ), .S0(quotient[2]), .Y(\u_div/PartRem[2][7] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_3_6  ( .A(\u_div/PartRem[4][6] ), .B(
        \u_div/SumTmp[3][6] ), .S0(quotient[3]), .Y(\u_div/PartRem[3][7] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_4_6  ( .A(\u_div/PartRem[5][6] ), .B(
        \u_div/SumTmp[4][6] ), .S0(quotient[4]), .Y(\u_div/PartRem[4][7] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_5_6  ( .A(\u_div/PartRem[6][6] ), .B(
        \u_div/SumTmp[5][6] ), .S0(quotient[5]), .Y(\u_div/PartRem[5][7] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_6_6  ( .A(\u_div/PartRem[7][6] ), .B(
        \u_div/SumTmp[6][6] ), .S0(quotient[6]), .Y(\u_div/PartRem[6][7] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_7_6  ( .A(\u_div/PartRem[8][6] ), .B(
        \u_div/SumTmp[7][6] ), .S0(quotient[7]), .Y(\u_div/PartRem[7][7] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_8_6  ( .A(\u_div/PartRem[9][6] ), .B(
        \u_div/SumTmp[8][6] ), .S0(quotient[8]), .Y(\u_div/PartRem[8][7] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_2_5  ( .A(\u_div/PartRem[3][5] ), .B(
        \u_div/SumTmp[2][5] ), .S0(quotient[2]), .Y(\u_div/PartRem[2][6] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_3_5  ( .A(\u_div/PartRem[4][5] ), .B(
        \u_div/SumTmp[3][5] ), .S0(quotient[3]), .Y(\u_div/PartRem[3][6] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_4_5  ( .A(\u_div/PartRem[5][5] ), .B(
        \u_div/SumTmp[4][5] ), .S0(quotient[4]), .Y(\u_div/PartRem[4][6] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_5_5  ( .A(\u_div/PartRem[6][5] ), .B(
        \u_div/SumTmp[5][5] ), .S0(quotient[5]), .Y(\u_div/PartRem[5][6] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_6_5  ( .A(\u_div/PartRem[7][5] ), .B(
        \u_div/SumTmp[6][5] ), .S0(quotient[6]), .Y(\u_div/PartRem[6][6] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_7_5  ( .A(\u_div/PartRem[8][5] ), .B(
        \u_div/SumTmp[7][5] ), .S0(quotient[7]), .Y(\u_div/PartRem[7][6] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_8_5  ( .A(\u_div/PartRem[9][5] ), .B(
        \u_div/SumTmp[8][5] ), .S0(quotient[8]), .Y(\u_div/PartRem[8][6] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_8_8  ( .A(\u_div/PartRem[9][8] ), .B(
        \u_div/SumTmp[8][8] ), .S0(quotient[8]), .Y(\u_div/PartRem[8][9] ) );
  MX2XL \u_div/u_mx_PartRem_0_1_5  ( .A(\u_div/PartRem[2][5] ), .B(
        \u_div/SumTmp[1][5] ), .S0(quotient[1]), .Y(\u_div/PartRem[1][6] ) );
  MX2XL \u_div/u_mx_PartRem_0_1_6  ( .A(\u_div/PartRem[2][6] ), .B(
        \u_div/SumTmp[1][6] ), .S0(quotient[1]), .Y(\u_div/PartRem[1][7] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_2_7  ( .A(\u_div/PartRem[3][7] ), .B(
        \u_div/SumTmp[2][7] ), .S0(quotient[2]), .Y(\u_div/PartRem[2][8] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_3_7  ( .A(\u_div/PartRem[4][7] ), .B(
        \u_div/SumTmp[3][7] ), .S0(quotient[3]), .Y(\u_div/PartRem[3][8] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_4_7  ( .A(\u_div/PartRem[5][7] ), .B(
        \u_div/SumTmp[4][7] ), .S0(quotient[4]), .Y(\u_div/PartRem[4][8] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_5_7  ( .A(\u_div/PartRem[6][7] ), .B(
        \u_div/SumTmp[5][7] ), .S0(quotient[5]), .Y(\u_div/PartRem[5][8] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_6_7  ( .A(\u_div/PartRem[7][7] ), .B(
        \u_div/SumTmp[6][7] ), .S0(quotient[6]), .Y(\u_div/PartRem[6][8] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_7_7  ( .A(\u_div/PartRem[8][7] ), .B(
        \u_div/SumTmp[7][7] ), .S0(quotient[7]), .Y(\u_div/PartRem[7][8] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_7_8  ( .A(\u_div/PartRem[8][8] ), .B(
        \u_div/SumTmp[7][8] ), .S0(quotient[7]), .Y(\u_div/PartRem[7][9] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_3_8  ( .A(\u_div/PartRem[4][8] ), .B(
        \u_div/SumTmp[3][8] ), .S0(quotient[3]), .Y(\u_div/PartRem[3][9] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_5_8  ( .A(\u_div/PartRem[6][8] ), .B(
        \u_div/SumTmp[5][8] ), .S0(quotient[5]), .Y(\u_div/PartRem[5][9] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_6_8  ( .A(\u_div/PartRem[7][8] ), .B(
        \u_div/SumTmp[6][8] ), .S0(quotient[6]), .Y(\u_div/PartRem[6][9] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_4_8  ( .A(\u_div/PartRem[5][8] ), .B(
        \u_div/SumTmp[4][8] ), .S0(quotient[4]), .Y(\u_div/PartRem[4][9] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_2_8  ( .A(\u_div/PartRem[3][8] ), .B(
        \u_div/SumTmp[2][8] ), .S0(quotient[2]), .Y(\u_div/PartRem[2][9] ) );
  OR2X2 U1 ( .A(\u_div/PartRem[2][9] ), .B(\u_div/u_add_PartRem_0_1/n2 ), .Y(
        quotient[1]) );
  MXI2XL U2 ( .A(\u_div/PartRem[2][3] ), .B(\u_div/SumTmp[1][3] ), .S0(
        quotient[1]), .Y(n1) );
  MXI2XL U3 ( .A(\u_div/SumTmp[1][2] ), .B(\u_div/SumTmp[1][2] ), .S0(
        quotient[1]), .Y(n2) );
  MXI2XL U4 ( .A(\u_div/PartRem[2][4] ), .B(\u_div/SumTmp[1][4] ), .S0(
        quotient[1]), .Y(n3) );
  CLKBUFX3 U5 ( .A(n35), .Y(quotient[3]) );
  OR2X1 U6 ( .A(\u_div/PartRem[4][9] ), .B(\u_div/u_add_PartRem_0_3/n2 ), .Y(
        n35) );
  CLKBUFX3 U7 ( .A(n33), .Y(quotient[5]) );
  OR2X1 U8 ( .A(\u_div/PartRem[6][9] ), .B(\u_div/u_add_PartRem_0_5/n2 ), .Y(
        n33) );
  CLKBUFX3 U9 ( .A(n34), .Y(quotient[4]) );
  OR2X1 U10 ( .A(\u_div/PartRem[5][9] ), .B(\u_div/u_add_PartRem_0_4/n2 ), .Y(
        n34) );
  CLKBUFX3 U11 ( .A(n36), .Y(quotient[2]) );
  OR2X1 U12 ( .A(\u_div/PartRem[3][9] ), .B(\u_div/u_add_PartRem_0_2/n2 ), .Y(
        n36) );
  CLKBUFX3 U13 ( .A(n32), .Y(quotient[6]) );
  OR2X1 U14 ( .A(\u_div/PartRem[7][9] ), .B(\u_div/u_add_PartRem_0_6/n2 ), .Y(
        n32) );
  CLKBUFX3 U15 ( .A(n31), .Y(quotient[7]) );
  OR2X1 U16 ( .A(\u_div/PartRem[8][9] ), .B(\u_div/u_add_PartRem_0_7/n2 ), .Y(
        n31) );
  CLKBUFX3 U17 ( .A(n30), .Y(quotient[8]) );
  OR2X1 U18 ( .A(\u_div/PartRem[9][9] ), .B(\u_div/u_add_PartRem_0_8/n2 ), .Y(
        n30) );
  NOR3X1 U19 ( .A(n1), .B(n2), .C(n3), .Y(n25) );
  CLKBUFX3 U20 ( .A(n27), .Y(n4) );
  CLKBUFX3 U21 ( .A(n29), .Y(n6) );
  OR2X1 U22 ( .A(\u_div/PartRem[10][9] ), .B(\u_div/u_add_PartRem_0_9/n2 ), 
        .Y(n29) );
  ADDHXL U23 ( .A(\u_div/SumTmp[19][0] ), .B(\u_div/u_add_PartRem_1_11/n2 ), 
        .CO(n27), .S(\u_div/SumTmp[11][8] ) );
  MXI2X1 U24 ( .A(\u_div/SumTmp[11][3] ), .B(\u_div/SumTmp[14][0] ), .S0(n4), 
        .Y(\u_div/PartRem[11][4] ) );
  CLKBUFX3 U25 ( .A(n28), .Y(n5) );
  OR2X1 U26 ( .A(\u_div/PartRem[11][9] ), .B(\u_div/u_add_PartRem_0_10/n2 ), 
        .Y(n28) );
  CLKINVX1 U27 ( .A(\u_div/SumTmp[14][0] ), .Y(\u_div/SumTmp[11][3] ) );
  XNOR2X1 U28 ( .A(\u_div/SumTmp[17][0] ), .B(\u_div/u_add_PartRem_1_11/n4 ), 
        .Y(\u_div/SumTmp[11][6] ) );
  NOR2X1 U29 ( .A(\u_div/u_add_PartRem_1_11/n4 ), .B(\u_div/SumTmp[17][0] ), 
        .Y(n14) );
  XOR2X1 U30 ( .A(\u_div/SumTmp[18][0] ), .B(n14), .Y(\u_div/SumTmp[11][7] )
         );
  NAND2BX1 U31 ( .AN(\u_div/SumTmp[18][0] ), .B(n14), .Y(
        \u_div/u_add_PartRem_1_11/n2 ) );
  CLKINVX1 U32 ( .A(\u_div/PartRem[11][3] ), .Y(\u_div/SumTmp[10][3] ) );
  XNOR2X1 U33 ( .A(\u_div/PartRem[11][6] ), .B(\u_div/u_add_PartRem_0_10/n5 ), 
        .Y(\u_div/SumTmp[10][6] ) );
  NOR2X1 U34 ( .A(\u_div/u_add_PartRem_0_10/n5 ), .B(\u_div/PartRem[11][6] ), 
        .Y(n15) );
  XOR2X1 U35 ( .A(\u_div/PartRem[11][7] ), .B(n15), .Y(\u_div/SumTmp[10][7] )
         );
  NAND2BX1 U36 ( .AN(\u_div/PartRem[11][7] ), .B(n15), .Y(
        \u_div/u_add_PartRem_0_10/n3 ) );
  CLKINVX1 U37 ( .A(\u_div/PartRem[10][3] ), .Y(\u_div/SumTmp[9][3] ) );
  XNOR2X1 U38 ( .A(\u_div/PartRem[10][6] ), .B(\u_div/u_add_PartRem_0_9/n5 ), 
        .Y(\u_div/SumTmp[9][6] ) );
  NOR2X1 U39 ( .A(\u_div/u_add_PartRem_0_9/n5 ), .B(\u_div/PartRem[10][6] ), 
        .Y(n16) );
  XOR2X1 U40 ( .A(\u_div/PartRem[10][7] ), .B(n16), .Y(\u_div/SumTmp[9][7] )
         );
  NAND2BX1 U41 ( .AN(\u_div/PartRem[10][7] ), .B(n16), .Y(
        \u_div/u_add_PartRem_0_9/n3 ) );
  CLKINVX1 U42 ( .A(\u_div/PartRem[9][3] ), .Y(\u_div/SumTmp[8][3] ) );
  XNOR2X1 U43 ( .A(\u_div/PartRem[9][6] ), .B(\u_div/u_add_PartRem_0_8/n5 ), 
        .Y(\u_div/SumTmp[8][6] ) );
  NOR2X1 U44 ( .A(\u_div/u_add_PartRem_0_8/n5 ), .B(\u_div/PartRem[9][6] ), 
        .Y(n17) );
  XOR2X1 U45 ( .A(\u_div/PartRem[9][7] ), .B(n17), .Y(\u_div/SumTmp[8][7] ) );
  NAND2BX1 U46 ( .AN(\u_div/PartRem[9][7] ), .B(n17), .Y(
        \u_div/u_add_PartRem_0_8/n3 ) );
  CLKINVX1 U47 ( .A(\u_div/PartRem[8][3] ), .Y(\u_div/SumTmp[7][3] ) );
  XNOR2X1 U48 ( .A(\u_div/PartRem[8][6] ), .B(\u_div/u_add_PartRem_0_7/n5 ), 
        .Y(\u_div/SumTmp[7][6] ) );
  NOR2X1 U49 ( .A(\u_div/u_add_PartRem_0_7/n5 ), .B(\u_div/PartRem[8][6] ), 
        .Y(n18) );
  XOR2X1 U50 ( .A(\u_div/PartRem[8][7] ), .B(n18), .Y(\u_div/SumTmp[7][7] ) );
  NAND2BX1 U51 ( .AN(\u_div/PartRem[8][7] ), .B(n18), .Y(
        \u_div/u_add_PartRem_0_7/n3 ) );
  CLKINVX1 U52 ( .A(\u_div/PartRem[7][3] ), .Y(\u_div/SumTmp[6][3] ) );
  XNOR2X1 U53 ( .A(\u_div/PartRem[7][6] ), .B(\u_div/u_add_PartRem_0_6/n5 ), 
        .Y(\u_div/SumTmp[6][6] ) );
  NOR2X1 U54 ( .A(\u_div/u_add_PartRem_0_6/n5 ), .B(\u_div/PartRem[7][6] ), 
        .Y(n19) );
  XOR2X1 U55 ( .A(\u_div/PartRem[7][7] ), .B(n19), .Y(\u_div/SumTmp[6][7] ) );
  NAND2BX1 U56 ( .AN(\u_div/PartRem[7][7] ), .B(n19), .Y(
        \u_div/u_add_PartRem_0_6/n3 ) );
  CLKINVX1 U57 ( .A(\u_div/PartRem[6][3] ), .Y(\u_div/SumTmp[5][3] ) );
  XNOR2X1 U58 ( .A(\u_div/PartRem[6][6] ), .B(\u_div/u_add_PartRem_0_5/n5 ), 
        .Y(\u_div/SumTmp[5][6] ) );
  NOR2X1 U59 ( .A(\u_div/u_add_PartRem_0_5/n5 ), .B(\u_div/PartRem[6][6] ), 
        .Y(n20) );
  XOR2X1 U60 ( .A(\u_div/PartRem[6][7] ), .B(n20), .Y(\u_div/SumTmp[5][7] ) );
  NAND2BX1 U61 ( .AN(\u_div/PartRem[6][7] ), .B(n20), .Y(
        \u_div/u_add_PartRem_0_5/n3 ) );
  CLKINVX1 U62 ( .A(\u_div/PartRem[5][3] ), .Y(\u_div/SumTmp[4][3] ) );
  XNOR2X1 U63 ( .A(\u_div/PartRem[5][6] ), .B(\u_div/u_add_PartRem_0_4/n5 ), 
        .Y(\u_div/SumTmp[4][6] ) );
  NOR2X1 U64 ( .A(\u_div/u_add_PartRem_0_4/n5 ), .B(\u_div/PartRem[5][6] ), 
        .Y(n21) );
  XOR2X1 U65 ( .A(\u_div/PartRem[5][7] ), .B(n21), .Y(\u_div/SumTmp[4][7] ) );
  NAND2BX1 U66 ( .AN(\u_div/PartRem[5][7] ), .B(n21), .Y(
        \u_div/u_add_PartRem_0_4/n3 ) );
  CLKINVX1 U67 ( .A(\u_div/PartRem[4][3] ), .Y(\u_div/SumTmp[3][3] ) );
  XNOR2X1 U68 ( .A(\u_div/PartRem[4][6] ), .B(\u_div/u_add_PartRem_0_3/n5 ), 
        .Y(\u_div/SumTmp[3][6] ) );
  NOR2X1 U69 ( .A(\u_div/u_add_PartRem_0_3/n5 ), .B(\u_div/PartRem[4][6] ), 
        .Y(n22) );
  XOR2X1 U70 ( .A(\u_div/PartRem[4][7] ), .B(n22), .Y(\u_div/SumTmp[3][7] ) );
  NAND2BX1 U71 ( .AN(\u_div/PartRem[4][7] ), .B(n22), .Y(
        \u_div/u_add_PartRem_0_3/n3 ) );
  CLKINVX1 U72 ( .A(\u_div/PartRem[3][3] ), .Y(\u_div/SumTmp[2][3] ) );
  XNOR2X1 U73 ( .A(\u_div/PartRem[3][6] ), .B(\u_div/u_add_PartRem_0_2/n5 ), 
        .Y(\u_div/SumTmp[2][6] ) );
  NOR2X1 U74 ( .A(\u_div/u_add_PartRem_0_2/n5 ), .B(\u_div/PartRem[3][6] ), 
        .Y(n23) );
  XOR2X1 U75 ( .A(\u_div/PartRem[3][7] ), .B(n23), .Y(\u_div/SumTmp[2][7] ) );
  NAND2BX1 U76 ( .AN(\u_div/PartRem[3][7] ), .B(n23), .Y(
        \u_div/u_add_PartRem_0_2/n3 ) );
  CLKINVX1 U77 ( .A(\u_div/PartRem[2][3] ), .Y(\u_div/SumTmp[1][3] ) );
  XNOR2X1 U78 ( .A(\u_div/PartRem[2][6] ), .B(\u_div/u_add_PartRem_0_1/n5 ), 
        .Y(\u_div/SumTmp[1][6] ) );
  NOR2X1 U79 ( .A(\u_div/u_add_PartRem_0_1/n5 ), .B(\u_div/PartRem[2][6] ), 
        .Y(n24) );
  XOR2X1 U80 ( .A(\u_div/PartRem[2][7] ), .B(n24), .Y(\u_div/SumTmp[1][7] ) );
  NAND2BX1 U81 ( .AN(\u_div/PartRem[2][7] ), .B(n24), .Y(
        \u_div/u_add_PartRem_0_1/n3 ) );
  OAI31XL U82 ( .A0(n25), .A1(\u_div/PartRem[1][7] ), .A2(
        \u_div/PartRem[1][6] ), .B0(\u_div/PartRem[1][8] ), .Y(n26) );
  NAND2BX1 U83 ( .AN(\u_div/PartRem[1][9] ), .B(n26), .Y(quotient[0]) );
endmodule


module CONT_DW01_add_33 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [19:1] carry;

  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  XOR3X1 U1_19 ( .A(A[19]), .B(B[19]), .C(carry[19]), .Y(SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  CMPR32X2 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  CMPR32X2 U1_16 ( .A(A[16]), .B(B[16]), .C(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  CMPR32X2 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module CONT_DW01_add_34 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [19:1] carry;

  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  XOR3X1 U1_19 ( .A(A[19]), .B(B[19]), .C(carry[19]), .Y(SUM[19]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2XL U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module CONT_DW_div_uns_11 ( a, b, quotient, remainder, divide_by_0 );
  input [19:0] a;
  input [8:0] b;
  output [19:0] quotient;
  output [8:0] remainder;
  output divide_by_0;
  wire   n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         \u_div/SumTmp[1][2] , \u_div/SumTmp[1][3] , \u_div/SumTmp[1][4] ,
         \u_div/SumTmp[1][5] , \u_div/SumTmp[1][6] , \u_div/SumTmp[1][7] ,
         \u_div/SumTmp[1][8] , \u_div/SumTmp[2][1] , \u_div/SumTmp[2][2] ,
         \u_div/SumTmp[2][3] , \u_div/SumTmp[2][4] , \u_div/SumTmp[2][5] ,
         \u_div/SumTmp[2][6] , \u_div/SumTmp[2][7] , \u_div/SumTmp[2][8] ,
         \u_div/SumTmp[3][0] , \u_div/SumTmp[3][1] , \u_div/SumTmp[3][2] ,
         \u_div/SumTmp[3][3] , \u_div/SumTmp[3][4] , \u_div/SumTmp[3][5] ,
         \u_div/SumTmp[3][6] , \u_div/SumTmp[3][7] , \u_div/SumTmp[3][8] ,
         \u_div/SumTmp[4][0] , \u_div/SumTmp[4][1] , \u_div/SumTmp[4][2] ,
         \u_div/SumTmp[4][3] , \u_div/SumTmp[4][4] , \u_div/SumTmp[4][5] ,
         \u_div/SumTmp[4][6] , \u_div/SumTmp[4][7] , \u_div/SumTmp[4][8] ,
         \u_div/SumTmp[5][0] , \u_div/SumTmp[5][1] , \u_div/SumTmp[5][2] ,
         \u_div/SumTmp[5][3] , \u_div/SumTmp[5][4] , \u_div/SumTmp[5][5] ,
         \u_div/SumTmp[5][6] , \u_div/SumTmp[5][7] , \u_div/SumTmp[5][8] ,
         \u_div/SumTmp[6][0] , \u_div/SumTmp[6][1] , \u_div/SumTmp[6][2] ,
         \u_div/SumTmp[6][3] , \u_div/SumTmp[6][4] , \u_div/SumTmp[6][5] ,
         \u_div/SumTmp[6][6] , \u_div/SumTmp[6][7] , \u_div/SumTmp[6][8] ,
         \u_div/SumTmp[7][0] , \u_div/SumTmp[7][1] , \u_div/SumTmp[7][2] ,
         \u_div/SumTmp[7][3] , \u_div/SumTmp[7][4] , \u_div/SumTmp[7][5] ,
         \u_div/SumTmp[7][6] , \u_div/SumTmp[7][7] , \u_div/SumTmp[7][8] ,
         \u_div/SumTmp[8][0] , \u_div/SumTmp[8][1] , \u_div/SumTmp[8][2] ,
         \u_div/SumTmp[8][3] , \u_div/SumTmp[8][4] , \u_div/SumTmp[8][5] ,
         \u_div/SumTmp[8][6] , \u_div/SumTmp[8][7] , \u_div/SumTmp[8][8] ,
         \u_div/SumTmp[9][0] , \u_div/SumTmp[9][1] , \u_div/SumTmp[9][2] ,
         \u_div/SumTmp[9][3] , \u_div/SumTmp[9][4] , \u_div/SumTmp[9][5] ,
         \u_div/SumTmp[9][6] , \u_div/SumTmp[9][7] , \u_div/SumTmp[9][8] ,
         \u_div/SumTmp[10][0] , \u_div/SumTmp[10][1] , \u_div/SumTmp[10][2] ,
         \u_div/SumTmp[10][3] , \u_div/SumTmp[10][4] , \u_div/SumTmp[10][5] ,
         \u_div/SumTmp[10][6] , \u_div/SumTmp[10][7] , \u_div/SumTmp[10][8] ,
         \u_div/SumTmp[11][0] , \u_div/SumTmp[11][1] , \u_div/SumTmp[11][2] ,
         \u_div/SumTmp[11][3] , \u_div/SumTmp[11][4] , \u_div/SumTmp[11][5] ,
         \u_div/SumTmp[11][6] , \u_div/SumTmp[11][7] , \u_div/SumTmp[11][8] ,
         \u_div/SumTmp[14][0] , \u_div/SumTmp[15][0] , \u_div/SumTmp[16][0] ,
         \u_div/SumTmp[17][0] , \u_div/SumTmp[18][0] , \u_div/SumTmp[19][0] ,
         \u_div/PartRem[1][6] , \u_div/PartRem[1][7] , \u_div/PartRem[1][8] ,
         \u_div/PartRem[1][9] , \u_div/PartRem[2][3] , \u_div/PartRem[2][4] ,
         \u_div/PartRem[2][5] , \u_div/PartRem[2][6] , \u_div/PartRem[2][7] ,
         \u_div/PartRem[2][8] , \u_div/PartRem[2][9] , \u_div/PartRem[3][3] ,
         \u_div/PartRem[3][4] , \u_div/PartRem[3][5] , \u_div/PartRem[3][6] ,
         \u_div/PartRem[3][7] , \u_div/PartRem[3][8] , \u_div/PartRem[3][9] ,
         \u_div/PartRem[4][3] , \u_div/PartRem[4][4] , \u_div/PartRem[4][5] ,
         \u_div/PartRem[4][6] , \u_div/PartRem[4][7] , \u_div/PartRem[4][8] ,
         \u_div/PartRem[4][9] , \u_div/PartRem[5][3] , \u_div/PartRem[5][4] ,
         \u_div/PartRem[5][5] , \u_div/PartRem[5][6] , \u_div/PartRem[5][7] ,
         \u_div/PartRem[5][8] , \u_div/PartRem[5][9] , \u_div/PartRem[6][3] ,
         \u_div/PartRem[6][4] , \u_div/PartRem[6][5] , \u_div/PartRem[6][6] ,
         \u_div/PartRem[6][7] , \u_div/PartRem[6][8] , \u_div/PartRem[6][9] ,
         \u_div/PartRem[7][3] , \u_div/PartRem[7][4] , \u_div/PartRem[7][5] ,
         \u_div/PartRem[7][6] , \u_div/PartRem[7][7] , \u_div/PartRem[7][8] ,
         \u_div/PartRem[7][9] , \u_div/PartRem[8][3] , \u_div/PartRem[8][4] ,
         \u_div/PartRem[8][5] , \u_div/PartRem[8][6] , \u_div/PartRem[8][7] ,
         \u_div/PartRem[8][8] , \u_div/PartRem[8][9] , \u_div/PartRem[9][3] ,
         \u_div/PartRem[9][4] , \u_div/PartRem[9][5] , \u_div/PartRem[9][6] ,
         \u_div/PartRem[9][7] , \u_div/PartRem[9][8] , \u_div/PartRem[9][9] ,
         \u_div/PartRem[10][3] , \u_div/PartRem[10][4] ,
         \u_div/PartRem[10][5] , \u_div/PartRem[10][6] ,
         \u_div/PartRem[10][7] , \u_div/PartRem[10][8] ,
         \u_div/PartRem[10][9] , \u_div/PartRem[11][3] ,
         \u_div/PartRem[11][4] , \u_div/PartRem[11][5] ,
         \u_div/PartRem[11][6] , \u_div/PartRem[11][7] ,
         \u_div/PartRem[11][8] , \u_div/PartRem[11][9] ,
         \u_div/u_add_PartRem_0_1/n6 , \u_div/u_add_PartRem_0_1/n5 ,
         \u_div/u_add_PartRem_0_1/n3 , \u_div/u_add_PartRem_0_1/n2 ,
         \u_div/u_add_PartRem_0_2/n6 , \u_div/u_add_PartRem_0_2/n5 ,
         \u_div/u_add_PartRem_0_2/n3 , \u_div/u_add_PartRem_0_2/n2 ,
         \u_div/u_add_PartRem_0_3/n6 , \u_div/u_add_PartRem_0_3/n5 ,
         \u_div/u_add_PartRem_0_3/n3 , \u_div/u_add_PartRem_0_3/n2 ,
         \u_div/u_add_PartRem_0_4/n6 , \u_div/u_add_PartRem_0_4/n5 ,
         \u_div/u_add_PartRem_0_4/n3 , \u_div/u_add_PartRem_0_4/n2 ,
         \u_div/u_add_PartRem_0_5/n6 , \u_div/u_add_PartRem_0_5/n5 ,
         \u_div/u_add_PartRem_0_5/n3 , \u_div/u_add_PartRem_0_5/n2 ,
         \u_div/u_add_PartRem_0_6/n6 , \u_div/u_add_PartRem_0_6/n5 ,
         \u_div/u_add_PartRem_0_6/n3 , \u_div/u_add_PartRem_0_6/n2 ,
         \u_div/u_add_PartRem_0_7/n6 , \u_div/u_add_PartRem_0_7/n5 ,
         \u_div/u_add_PartRem_0_7/n3 , \u_div/u_add_PartRem_0_7/n2 ,
         \u_div/u_add_PartRem_0_8/n6 , \u_div/u_add_PartRem_0_8/n5 ,
         \u_div/u_add_PartRem_0_8/n3 , \u_div/u_add_PartRem_0_8/n2 ,
         \u_div/u_add_PartRem_0_9/n6 , \u_div/u_add_PartRem_0_9/n5 ,
         \u_div/u_add_PartRem_0_9/n3 , \u_div/u_add_PartRem_0_9/n2 ,
         \u_div/u_add_PartRem_0_10/n6 , \u_div/u_add_PartRem_0_10/n5 ,
         \u_div/u_add_PartRem_0_10/n3 , \u_div/u_add_PartRem_0_10/n2 ,
         \u_div/u_add_PartRem_1_11/n5 , \u_div/u_add_PartRem_1_11/n4 ,
         \u_div/u_add_PartRem_1_11/n2 , n1, n2, n3, n4, n5, n6, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign \u_div/SumTmp[3][0]  = a[3];
  assign \u_div/SumTmp[4][0]  = a[4];
  assign \u_div/SumTmp[5][0]  = a[5];
  assign \u_div/SumTmp[6][0]  = a[6];
  assign \u_div/SumTmp[7][0]  = a[7];
  assign \u_div/SumTmp[8][0]  = a[8];
  assign \u_div/SumTmp[9][0]  = a[9];
  assign \u_div/SumTmp[10][0]  = a[10];
  assign \u_div/SumTmp[11][0]  = a[11];
  assign \u_div/SumTmp[11][1]  = a[12];
  assign \u_div/SumTmp[11][2]  = a[13];
  assign \u_div/SumTmp[14][0]  = a[14];
  assign \u_div/SumTmp[15][0]  = a[15];
  assign \u_div/SumTmp[16][0]  = a[16];
  assign \u_div/SumTmp[17][0]  = a[17];
  assign \u_div/SumTmp[18][0]  = a[18];
  assign \u_div/SumTmp[19][0]  = a[19];

  ADDHXL \u_div/u_add_PartRem_0_1/U9  ( .A(\u_div/PartRem[2][4] ), .B(
        \u_div/PartRem[2][3] ), .CO(\u_div/u_add_PartRem_0_1/n6 ), .S(
        \u_div/SumTmp[1][4] ) );
  ADDHXL \u_div/u_add_PartRem_0_1/U8  ( .A(\u_div/PartRem[2][5] ), .B(
        \u_div/u_add_PartRem_0_1/n6 ), .CO(\u_div/u_add_PartRem_0_1/n5 ), .S(
        \u_div/SumTmp[1][5] ) );
  ADDHXL \u_div/u_add_PartRem_0_1/U3  ( .A(\u_div/PartRem[2][8] ), .B(
        \u_div/u_add_PartRem_0_1/n3 ), .CO(\u_div/u_add_PartRem_0_1/n2 ), .S(
        \u_div/SumTmp[1][8] ) );
  ADDHXL \u_div/u_add_PartRem_0_2/U9  ( .A(\u_div/PartRem[3][4] ), .B(
        \u_div/PartRem[3][3] ), .CO(\u_div/u_add_PartRem_0_2/n6 ), .S(
        \u_div/SumTmp[2][4] ) );
  ADDHXL \u_div/u_add_PartRem_0_2/U8  ( .A(\u_div/PartRem[3][5] ), .B(
        \u_div/u_add_PartRem_0_2/n6 ), .CO(\u_div/u_add_PartRem_0_2/n5 ), .S(
        \u_div/SumTmp[2][5] ) );
  ADDHXL \u_div/u_add_PartRem_0_2/U3  ( .A(\u_div/PartRem[3][8] ), .B(
        \u_div/u_add_PartRem_0_2/n3 ), .CO(\u_div/u_add_PartRem_0_2/n2 ), .S(
        \u_div/SumTmp[2][8] ) );
  ADDHXL \u_div/u_add_PartRem_0_3/U9  ( .A(\u_div/PartRem[4][4] ), .B(
        \u_div/PartRem[4][3] ), .CO(\u_div/u_add_PartRem_0_3/n6 ), .S(
        \u_div/SumTmp[3][4] ) );
  ADDHXL \u_div/u_add_PartRem_0_3/U8  ( .A(\u_div/PartRem[4][5] ), .B(
        \u_div/u_add_PartRem_0_3/n6 ), .CO(\u_div/u_add_PartRem_0_3/n5 ), .S(
        \u_div/SumTmp[3][5] ) );
  ADDHXL \u_div/u_add_PartRem_0_3/U3  ( .A(\u_div/PartRem[4][8] ), .B(
        \u_div/u_add_PartRem_0_3/n3 ), .CO(\u_div/u_add_PartRem_0_3/n2 ), .S(
        \u_div/SumTmp[3][8] ) );
  ADDHXL \u_div/u_add_PartRem_0_4/U9  ( .A(\u_div/PartRem[5][4] ), .B(
        \u_div/PartRem[5][3] ), .CO(\u_div/u_add_PartRem_0_4/n6 ), .S(
        \u_div/SumTmp[4][4] ) );
  ADDHXL \u_div/u_add_PartRem_0_4/U8  ( .A(\u_div/PartRem[5][5] ), .B(
        \u_div/u_add_PartRem_0_4/n6 ), .CO(\u_div/u_add_PartRem_0_4/n5 ), .S(
        \u_div/SumTmp[4][5] ) );
  ADDHXL \u_div/u_add_PartRem_0_4/U3  ( .A(\u_div/PartRem[5][8] ), .B(
        \u_div/u_add_PartRem_0_4/n3 ), .CO(\u_div/u_add_PartRem_0_4/n2 ), .S(
        \u_div/SumTmp[4][8] ) );
  ADDHXL \u_div/u_add_PartRem_0_5/U9  ( .A(\u_div/PartRem[6][4] ), .B(
        \u_div/PartRem[6][3] ), .CO(\u_div/u_add_PartRem_0_5/n6 ), .S(
        \u_div/SumTmp[5][4] ) );
  ADDHXL \u_div/u_add_PartRem_0_5/U8  ( .A(\u_div/PartRem[6][5] ), .B(
        \u_div/u_add_PartRem_0_5/n6 ), .CO(\u_div/u_add_PartRem_0_5/n5 ), .S(
        \u_div/SumTmp[5][5] ) );
  ADDHXL \u_div/u_add_PartRem_0_5/U3  ( .A(\u_div/PartRem[6][8] ), .B(
        \u_div/u_add_PartRem_0_5/n3 ), .CO(\u_div/u_add_PartRem_0_5/n2 ), .S(
        \u_div/SumTmp[5][8] ) );
  ADDHXL \u_div/u_add_PartRem_0_6/U9  ( .A(\u_div/PartRem[7][4] ), .B(
        \u_div/PartRem[7][3] ), .CO(\u_div/u_add_PartRem_0_6/n6 ), .S(
        \u_div/SumTmp[6][4] ) );
  ADDHXL \u_div/u_add_PartRem_0_6/U8  ( .A(\u_div/PartRem[7][5] ), .B(
        \u_div/u_add_PartRem_0_6/n6 ), .CO(\u_div/u_add_PartRem_0_6/n5 ), .S(
        \u_div/SumTmp[6][5] ) );
  ADDHXL \u_div/u_add_PartRem_0_6/U3  ( .A(\u_div/PartRem[7][8] ), .B(
        \u_div/u_add_PartRem_0_6/n3 ), .CO(\u_div/u_add_PartRem_0_6/n2 ), .S(
        \u_div/SumTmp[6][8] ) );
  ADDHXL \u_div/u_add_PartRem_0_7/U9  ( .A(\u_div/PartRem[8][4] ), .B(
        \u_div/PartRem[8][3] ), .CO(\u_div/u_add_PartRem_0_7/n6 ), .S(
        \u_div/SumTmp[7][4] ) );
  ADDHXL \u_div/u_add_PartRem_0_7/U8  ( .A(\u_div/PartRem[8][5] ), .B(
        \u_div/u_add_PartRem_0_7/n6 ), .CO(\u_div/u_add_PartRem_0_7/n5 ), .S(
        \u_div/SumTmp[7][5] ) );
  ADDHXL \u_div/u_add_PartRem_0_7/U3  ( .A(\u_div/PartRem[8][8] ), .B(
        \u_div/u_add_PartRem_0_7/n3 ), .CO(\u_div/u_add_PartRem_0_7/n2 ), .S(
        \u_div/SumTmp[7][8] ) );
  ADDHXL \u_div/u_add_PartRem_0_8/U9  ( .A(\u_div/PartRem[9][4] ), .B(
        \u_div/PartRem[9][3] ), .CO(\u_div/u_add_PartRem_0_8/n6 ), .S(
        \u_div/SumTmp[8][4] ) );
  ADDHXL \u_div/u_add_PartRem_0_8/U8  ( .A(\u_div/PartRem[9][5] ), .B(
        \u_div/u_add_PartRem_0_8/n6 ), .CO(\u_div/u_add_PartRem_0_8/n5 ), .S(
        \u_div/SumTmp[8][5] ) );
  ADDHXL \u_div/u_add_PartRem_0_8/U3  ( .A(\u_div/PartRem[9][8] ), .B(
        \u_div/u_add_PartRem_0_8/n3 ), .CO(\u_div/u_add_PartRem_0_8/n2 ), .S(
        \u_div/SumTmp[8][8] ) );
  ADDHXL \u_div/u_add_PartRem_0_9/U9  ( .A(\u_div/PartRem[10][4] ), .B(
        \u_div/PartRem[10][3] ), .CO(\u_div/u_add_PartRem_0_9/n6 ), .S(
        \u_div/SumTmp[9][4] ) );
  ADDHXL \u_div/u_add_PartRem_0_9/U8  ( .A(\u_div/PartRem[10][5] ), .B(
        \u_div/u_add_PartRem_0_9/n6 ), .CO(\u_div/u_add_PartRem_0_9/n5 ), .S(
        \u_div/SumTmp[9][5] ) );
  ADDHXL \u_div/u_add_PartRem_0_9/U3  ( .A(\u_div/PartRem[10][8] ), .B(
        \u_div/u_add_PartRem_0_9/n3 ), .CO(\u_div/u_add_PartRem_0_9/n2 ), .S(
        \u_div/SumTmp[9][8] ) );
  ADDHXL \u_div/u_add_PartRem_0_10/U9  ( .A(\u_div/PartRem[11][4] ), .B(
        \u_div/PartRem[11][3] ), .CO(\u_div/u_add_PartRem_0_10/n6 ), .S(
        \u_div/SumTmp[10][4] ) );
  ADDHXL \u_div/u_add_PartRem_0_10/U8  ( .A(\u_div/PartRem[11][5] ), .B(
        \u_div/u_add_PartRem_0_10/n6 ), .CO(\u_div/u_add_PartRem_0_10/n5 ), 
        .S(\u_div/SumTmp[10][5] ) );
  ADDHXL \u_div/u_add_PartRem_0_10/U3  ( .A(\u_div/PartRem[11][8] ), .B(
        \u_div/u_add_PartRem_0_10/n3 ), .CO(\u_div/u_add_PartRem_0_10/n2 ), 
        .S(\u_div/SumTmp[10][8] ) );
  ADDHXL \u_div/u_add_PartRem_1_11/U8  ( .A(\u_div/SumTmp[15][0] ), .B(
        \u_div/SumTmp[14][0] ), .CO(\u_div/u_add_PartRem_1_11/n5 ), .S(
        \u_div/SumTmp[11][4] ) );
  ADDHXL \u_div/u_add_PartRem_1_11/U7  ( .A(\u_div/SumTmp[16][0] ), .B(
        \u_div/u_add_PartRem_1_11/n5 ), .CO(\u_div/u_add_PartRem_1_11/n4 ), 
        .S(\u_div/SumTmp[11][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_3_0  ( .A(\u_div/SumTmp[3][0] ), .B(
        \u_div/SumTmp[3][0] ), .S0(quotient[3]), .Y(\u_div/SumTmp[2][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_2_1  ( .A(\u_div/SumTmp[2][1] ), .B(
        \u_div/SumTmp[2][1] ), .S0(quotient[2]), .Y(\u_div/SumTmp[1][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_11_7  ( .A(\u_div/SumTmp[18][0] ), .B(
        \u_div/SumTmp[11][7] ), .S0(n4), .Y(\u_div/PartRem[11][8] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_11_6  ( .A(\u_div/SumTmp[17][0] ), .B(
        \u_div/SumTmp[11][6] ), .S0(n4), .Y(\u_div/PartRem[11][7] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_11_8  ( .A(\u_div/SumTmp[19][0] ), .B(
        \u_div/SumTmp[11][8] ), .S0(n4), .Y(\u_div/PartRem[11][9] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_11_3  ( .A(\u_div/SumTmp[14][0] ), .B(
        \u_div/SumTmp[11][3] ), .S0(n4), .Y(\u_div/PartRem[11][4] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_11_4  ( .A(\u_div/SumTmp[15][0] ), .B(
        \u_div/SumTmp[11][4] ), .S0(n4), .Y(\u_div/PartRem[11][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_5_0  ( .A(\u_div/SumTmp[5][0] ), .B(
        \u_div/SumTmp[5][0] ), .S0(quotient[5]), .Y(\u_div/SumTmp[4][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_4_1  ( .A(\u_div/SumTmp[4][1] ), .B(
        \u_div/SumTmp[4][1] ), .S0(quotient[4]), .Y(\u_div/SumTmp[3][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_3_2  ( .A(\u_div/SumTmp[3][2] ), .B(
        \u_div/SumTmp[3][2] ), .S0(quotient[3]), .Y(\u_div/PartRem[3][3] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_6_0  ( .A(\u_div/SumTmp[6][0] ), .B(
        \u_div/SumTmp[6][0] ), .S0(quotient[6]), .Y(\u_div/SumTmp[5][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_5_1  ( .A(\u_div/SumTmp[5][1] ), .B(
        \u_div/SumTmp[5][1] ), .S0(quotient[5]), .Y(\u_div/SumTmp[4][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_4_2  ( .A(\u_div/SumTmp[4][2] ), .B(
        \u_div/SumTmp[4][2] ), .S0(quotient[4]), .Y(\u_div/PartRem[4][3] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_7_0  ( .A(\u_div/SumTmp[7][0] ), .B(
        \u_div/SumTmp[7][0] ), .S0(quotient[7]), .Y(\u_div/SumTmp[6][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_6_1  ( .A(\u_div/SumTmp[6][1] ), .B(
        \u_div/SumTmp[6][1] ), .S0(quotient[6]), .Y(\u_div/SumTmp[5][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_5_2  ( .A(\u_div/SumTmp[5][2] ), .B(
        \u_div/SumTmp[5][2] ), .S0(quotient[5]), .Y(\u_div/PartRem[5][3] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_8_0  ( .A(\u_div/SumTmp[8][0] ), .B(
        \u_div/SumTmp[8][0] ), .S0(quotient[8]), .Y(\u_div/SumTmp[7][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_7_1  ( .A(\u_div/SumTmp[7][1] ), .B(
        \u_div/SumTmp[7][1] ), .S0(quotient[7]), .Y(\u_div/SumTmp[6][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_6_2  ( .A(\u_div/SumTmp[6][2] ), .B(
        \u_div/SumTmp[6][2] ), .S0(quotient[6]), .Y(\u_div/PartRem[6][3] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_9_0  ( .A(\u_div/SumTmp[9][0] ), .B(
        \u_div/SumTmp[9][0] ), .S0(n6), .Y(\u_div/SumTmp[8][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_8_1  ( .A(\u_div/SumTmp[8][1] ), .B(
        \u_div/SumTmp[8][1] ), .S0(quotient[8]), .Y(\u_div/SumTmp[7][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_7_2  ( .A(\u_div/SumTmp[7][2] ), .B(
        \u_div/SumTmp[7][2] ), .S0(quotient[7]), .Y(\u_div/PartRem[7][3] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_10_0  ( .A(\u_div/SumTmp[10][0] ), .B(
        \u_div/SumTmp[10][0] ), .S0(n5), .Y(\u_div/SumTmp[9][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_9_1  ( .A(\u_div/SumTmp[9][1] ), .B(
        \u_div/SumTmp[9][1] ), .S0(n6), .Y(\u_div/SumTmp[8][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_8_2  ( .A(\u_div/SumTmp[8][2] ), .B(
        \u_div/SumTmp[8][2] ), .S0(quotient[8]), .Y(\u_div/PartRem[8][3] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_4_0  ( .A(\u_div/SumTmp[4][0] ), .B(
        \u_div/SumTmp[4][0] ), .S0(quotient[4]), .Y(\u_div/SumTmp[3][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_3_1  ( .A(\u_div/SumTmp[3][1] ), .B(
        \u_div/SumTmp[3][1] ), .S0(quotient[3]), .Y(\u_div/SumTmp[2][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_2_2  ( .A(\u_div/SumTmp[2][2] ), .B(
        \u_div/SumTmp[2][2] ), .S0(quotient[2]), .Y(\u_div/PartRem[2][3] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_11_0  ( .A(\u_div/SumTmp[11][0] ), .B(
        \u_div/SumTmp[11][0] ), .S0(n4), .Y(\u_div/SumTmp[10][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_10_1  ( .A(\u_div/SumTmp[10][1] ), .B(
        \u_div/SumTmp[10][1] ), .S0(n5), .Y(\u_div/SumTmp[9][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_9_2  ( .A(\u_div/SumTmp[9][2] ), .B(
        \u_div/SumTmp[9][2] ), .S0(n6), .Y(\u_div/PartRem[9][3] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_11_1  ( .A(\u_div/SumTmp[11][1] ), .B(
        \u_div/SumTmp[11][1] ), .S0(n4), .Y(\u_div/SumTmp[10][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_10_2  ( .A(\u_div/SumTmp[10][2] ), .B(
        \u_div/SumTmp[10][2] ), .S0(n5), .Y(\u_div/PartRem[10][3] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_11_2  ( .A(\u_div/SumTmp[11][2] ), .B(
        \u_div/SumTmp[11][2] ), .S0(n4), .Y(\u_div/PartRem[11][3] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_11_5  ( .A(\u_div/SumTmp[16][0] ), .B(
        \u_div/SumTmp[11][5] ), .S0(n4), .Y(\u_div/PartRem[11][6] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_10_7  ( .A(\u_div/PartRem[11][7] ), .B(
        \u_div/SumTmp[10][7] ), .S0(n5), .Y(\u_div/PartRem[10][8] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_10_6  ( .A(\u_div/PartRem[11][6] ), .B(
        \u_div/SumTmp[10][6] ), .S0(n5), .Y(\u_div/PartRem[10][7] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_10_8  ( .A(\u_div/PartRem[11][8] ), .B(
        \u_div/SumTmp[10][8] ), .S0(n5), .Y(\u_div/PartRem[10][9] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_3_3  ( .A(\u_div/PartRem[4][3] ), .B(
        \u_div/SumTmp[3][3] ), .S0(quotient[3]), .Y(\u_div/PartRem[3][4] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_4_3  ( .A(\u_div/PartRem[5][3] ), .B(
        \u_div/SumTmp[4][3] ), .S0(quotient[4]), .Y(\u_div/PartRem[4][4] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_5_3  ( .A(\u_div/PartRem[6][3] ), .B(
        \u_div/SumTmp[5][3] ), .S0(quotient[5]), .Y(\u_div/PartRem[5][4] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_6_3  ( .A(\u_div/PartRem[7][3] ), .B(
        \u_div/SumTmp[6][3] ), .S0(quotient[6]), .Y(\u_div/PartRem[6][4] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_7_3  ( .A(\u_div/PartRem[8][3] ), .B(
        \u_div/SumTmp[7][3] ), .S0(quotient[7]), .Y(\u_div/PartRem[7][4] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_8_3  ( .A(\u_div/PartRem[9][3] ), .B(
        \u_div/SumTmp[8][3] ), .S0(quotient[8]), .Y(\u_div/PartRem[8][4] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_2_3  ( .A(\u_div/PartRem[3][3] ), .B(
        \u_div/SumTmp[2][3] ), .S0(quotient[2]), .Y(\u_div/PartRem[2][4] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_9_3  ( .A(\u_div/PartRem[10][3] ), .B(
        \u_div/SumTmp[9][3] ), .S0(n6), .Y(\u_div/PartRem[9][4] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_10_3  ( .A(\u_div/PartRem[11][3] ), .B(
        \u_div/SumTmp[10][3] ), .S0(n5), .Y(\u_div/PartRem[10][4] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_10_4  ( .A(\u_div/PartRem[11][4] ), .B(
        \u_div/SumTmp[10][4] ), .S0(n5), .Y(\u_div/PartRem[10][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_10_5  ( .A(\u_div/PartRem[11][5] ), .B(
        \u_div/SumTmp[10][5] ), .S0(n5), .Y(\u_div/PartRem[10][6] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_9_7  ( .A(\u_div/PartRem[10][7] ), .B(
        \u_div/SumTmp[9][7] ), .S0(n6), .Y(\u_div/PartRem[9][8] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_9_6  ( .A(\u_div/PartRem[10][6] ), .B(
        \u_div/SumTmp[9][6] ), .S0(n6), .Y(\u_div/PartRem[9][7] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_9_8  ( .A(\u_div/PartRem[10][8] ), .B(
        \u_div/SumTmp[9][8] ), .S0(n6), .Y(\u_div/PartRem[9][9] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_2_4  ( .A(\u_div/PartRem[3][4] ), .B(
        \u_div/SumTmp[2][4] ), .S0(quotient[2]), .Y(\u_div/PartRem[2][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_3_4  ( .A(\u_div/PartRem[4][4] ), .B(
        \u_div/SumTmp[3][4] ), .S0(quotient[3]), .Y(\u_div/PartRem[3][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_4_4  ( .A(\u_div/PartRem[5][4] ), .B(
        \u_div/SumTmp[4][4] ), .S0(quotient[4]), .Y(\u_div/PartRem[4][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_5_4  ( .A(\u_div/PartRem[6][4] ), .B(
        \u_div/SumTmp[5][4] ), .S0(quotient[5]), .Y(\u_div/PartRem[5][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_6_4  ( .A(\u_div/PartRem[7][4] ), .B(
        \u_div/SumTmp[6][4] ), .S0(quotient[6]), .Y(\u_div/PartRem[6][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_7_4  ( .A(\u_div/PartRem[8][4] ), .B(
        \u_div/SumTmp[7][4] ), .S0(quotient[7]), .Y(\u_div/PartRem[7][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_8_4  ( .A(\u_div/PartRem[9][4] ), .B(
        \u_div/SumTmp[8][4] ), .S0(quotient[8]), .Y(\u_div/PartRem[8][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_9_4  ( .A(\u_div/PartRem[10][4] ), .B(
        \u_div/SumTmp[9][4] ), .S0(n6), .Y(\u_div/PartRem[9][5] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_9_5  ( .A(\u_div/PartRem[10][5] ), .B(
        \u_div/SumTmp[9][5] ), .S0(n6), .Y(\u_div/PartRem[9][6] ) );
  MX2XL \u_div/u_mx_PartRem_0_1_7  ( .A(\u_div/PartRem[2][7] ), .B(
        \u_div/SumTmp[1][7] ), .S0(quotient[1]), .Y(\u_div/PartRem[1][8] ) );
  MX2XL \u_div/u_mx_PartRem_0_1_8  ( .A(\u_div/PartRem[2][8] ), .B(
        \u_div/SumTmp[1][8] ), .S0(quotient[1]), .Y(\u_div/PartRem[1][9] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_8_7  ( .A(\u_div/PartRem[9][7] ), .B(
        \u_div/SumTmp[8][7] ), .S0(quotient[8]), .Y(\u_div/PartRem[8][8] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_2_6  ( .A(\u_div/PartRem[3][6] ), .B(
        \u_div/SumTmp[2][6] ), .S0(quotient[2]), .Y(\u_div/PartRem[2][7] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_3_6  ( .A(\u_div/PartRem[4][6] ), .B(
        \u_div/SumTmp[3][6] ), .S0(quotient[3]), .Y(\u_div/PartRem[3][7] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_4_6  ( .A(\u_div/PartRem[5][6] ), .B(
        \u_div/SumTmp[4][6] ), .S0(quotient[4]), .Y(\u_div/PartRem[4][7] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_5_6  ( .A(\u_div/PartRem[6][6] ), .B(
        \u_div/SumTmp[5][6] ), .S0(quotient[5]), .Y(\u_div/PartRem[5][7] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_6_6  ( .A(\u_div/PartRem[7][6] ), .B(
        \u_div/SumTmp[6][6] ), .S0(quotient[6]), .Y(\u_div/PartRem[6][7] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_7_6  ( .A(\u_div/PartRem[8][6] ), .B(
        \u_div/SumTmp[7][6] ), .S0(quotient[7]), .Y(\u_div/PartRem[7][7] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_8_6  ( .A(\u_div/PartRem[9][6] ), .B(
        \u_div/SumTmp[8][6] ), .S0(quotient[8]), .Y(\u_div/PartRem[8][7] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_2_5  ( .A(\u_div/PartRem[3][5] ), .B(
        \u_div/SumTmp[2][5] ), .S0(quotient[2]), .Y(\u_div/PartRem[2][6] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_8_8  ( .A(\u_div/PartRem[9][8] ), .B(
        \u_div/SumTmp[8][8] ), .S0(quotient[8]), .Y(\u_div/PartRem[8][9] ) );
  MX2XL \u_div/u_mx_PartRem_0_1_5  ( .A(\u_div/PartRem[2][5] ), .B(
        \u_div/SumTmp[1][5] ), .S0(quotient[1]), .Y(\u_div/PartRem[1][6] ) );
  MX2XL \u_div/u_mx_PartRem_0_1_6  ( .A(\u_div/PartRem[2][6] ), .B(
        \u_div/SumTmp[1][6] ), .S0(quotient[1]), .Y(\u_div/PartRem[1][7] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_3_5  ( .A(\u_div/PartRem[4][5] ), .B(
        \u_div/SumTmp[3][5] ), .S0(quotient[3]), .Y(\u_div/PartRem[3][6] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_4_5  ( .A(\u_div/PartRem[5][5] ), .B(
        \u_div/SumTmp[4][5] ), .S0(quotient[4]), .Y(\u_div/PartRem[4][6] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_5_5  ( .A(\u_div/PartRem[6][5] ), .B(
        \u_div/SumTmp[5][5] ), .S0(quotient[5]), .Y(\u_div/PartRem[5][6] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_6_5  ( .A(\u_div/PartRem[7][5] ), .B(
        \u_div/SumTmp[6][5] ), .S0(quotient[6]), .Y(\u_div/PartRem[6][6] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_7_5  ( .A(\u_div/PartRem[8][5] ), .B(
        \u_div/SumTmp[7][5] ), .S0(quotient[7]), .Y(\u_div/PartRem[7][6] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_8_5  ( .A(\u_div/PartRem[9][5] ), .B(
        \u_div/SumTmp[8][5] ), .S0(quotient[8]), .Y(\u_div/PartRem[8][6] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_2_7  ( .A(\u_div/PartRem[3][7] ), .B(
        \u_div/SumTmp[2][7] ), .S0(quotient[2]), .Y(\u_div/PartRem[2][8] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_3_7  ( .A(\u_div/PartRem[4][7] ), .B(
        \u_div/SumTmp[3][7] ), .S0(quotient[3]), .Y(\u_div/PartRem[3][8] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_4_7  ( .A(\u_div/PartRem[5][7] ), .B(
        \u_div/SumTmp[4][7] ), .S0(quotient[4]), .Y(\u_div/PartRem[4][8] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_5_7  ( .A(\u_div/PartRem[6][7] ), .B(
        \u_div/SumTmp[5][7] ), .S0(quotient[5]), .Y(\u_div/PartRem[5][8] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_6_7  ( .A(\u_div/PartRem[7][7] ), .B(
        \u_div/SumTmp[6][7] ), .S0(quotient[6]), .Y(\u_div/PartRem[6][8] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_7_7  ( .A(\u_div/PartRem[8][7] ), .B(
        \u_div/SumTmp[7][7] ), .S0(quotient[7]), .Y(\u_div/PartRem[7][8] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_7_8  ( .A(\u_div/PartRem[8][8] ), .B(
        \u_div/SumTmp[7][8] ), .S0(quotient[7]), .Y(\u_div/PartRem[7][9] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_5_8  ( .A(\u_div/PartRem[6][8] ), .B(
        \u_div/SumTmp[5][8] ), .S0(quotient[5]), .Y(\u_div/PartRem[5][9] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_3_8  ( .A(\u_div/PartRem[4][8] ), .B(
        \u_div/SumTmp[3][8] ), .S0(quotient[3]), .Y(\u_div/PartRem[3][9] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_4_8  ( .A(\u_div/PartRem[5][8] ), .B(
        \u_div/SumTmp[4][8] ), .S0(quotient[4]), .Y(\u_div/PartRem[4][9] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_6_8  ( .A(\u_div/PartRem[7][8] ), .B(
        \u_div/SumTmp[6][8] ), .S0(quotient[6]), .Y(\u_div/PartRem[6][9] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_2_8  ( .A(\u_div/PartRem[3][8] ), .B(
        \u_div/SumTmp[2][8] ), .S0(quotient[2]), .Y(\u_div/PartRem[2][9] ) );
  OR2X2 U1 ( .A(\u_div/PartRem[2][9] ), .B(\u_div/u_add_PartRem_0_1/n2 ), .Y(
        quotient[1]) );
  MXI2XL U2 ( .A(\u_div/PartRem[2][3] ), .B(\u_div/SumTmp[1][3] ), .S0(
        quotient[1]), .Y(n1) );
  MXI2XL U3 ( .A(\u_div/SumTmp[1][2] ), .B(\u_div/SumTmp[1][2] ), .S0(
        quotient[1]), .Y(n2) );
  MXI2XL U4 ( .A(\u_div/PartRem[2][4] ), .B(\u_div/SumTmp[1][4] ), .S0(
        quotient[1]), .Y(n3) );
  CLKBUFX3 U5 ( .A(n33), .Y(quotient[5]) );
  OR2X1 U6 ( .A(\u_div/PartRem[6][9] ), .B(\u_div/u_add_PartRem_0_5/n2 ), .Y(
        n33) );
  CLKBUFX3 U7 ( .A(n35), .Y(quotient[3]) );
  OR2X1 U8 ( .A(\u_div/PartRem[4][9] ), .B(\u_div/u_add_PartRem_0_3/n2 ), .Y(
        n35) );
  CLKBUFX3 U9 ( .A(n36), .Y(quotient[2]) );
  OR2X1 U10 ( .A(\u_div/PartRem[3][9] ), .B(\u_div/u_add_PartRem_0_2/n2 ), .Y(
        n36) );
  CLKBUFX3 U11 ( .A(n34), .Y(quotient[4]) );
  OR2X1 U12 ( .A(\u_div/PartRem[5][9] ), .B(\u_div/u_add_PartRem_0_4/n2 ), .Y(
        n34) );
  CLKBUFX3 U13 ( .A(n32), .Y(quotient[6]) );
  OR2X1 U14 ( .A(\u_div/PartRem[7][9] ), .B(\u_div/u_add_PartRem_0_6/n2 ), .Y(
        n32) );
  CLKBUFX3 U15 ( .A(n31), .Y(quotient[7]) );
  OR2X1 U16 ( .A(\u_div/PartRem[8][9] ), .B(\u_div/u_add_PartRem_0_7/n2 ), .Y(
        n31) );
  CLKBUFX3 U17 ( .A(n30), .Y(quotient[8]) );
  OR2X1 U18 ( .A(\u_div/PartRem[9][9] ), .B(\u_div/u_add_PartRem_0_8/n2 ), .Y(
        n30) );
  NOR3X1 U19 ( .A(n1), .B(n2), .C(n3), .Y(n25) );
  CLKBUFX3 U20 ( .A(n27), .Y(n4) );
  CLKBUFX3 U21 ( .A(n29), .Y(n6) );
  OR2X1 U22 ( .A(\u_div/PartRem[10][9] ), .B(\u_div/u_add_PartRem_0_9/n2 ), 
        .Y(n29) );
  ADDHXL U23 ( .A(\u_div/SumTmp[19][0] ), .B(\u_div/u_add_PartRem_1_11/n2 ), 
        .CO(n27), .S(\u_div/SumTmp[11][8] ) );
  CLKBUFX3 U24 ( .A(n28), .Y(n5) );
  OR2X1 U25 ( .A(\u_div/PartRem[11][9] ), .B(\u_div/u_add_PartRem_0_10/n2 ), 
        .Y(n28) );
  CLKINVX1 U26 ( .A(\u_div/SumTmp[14][0] ), .Y(\u_div/SumTmp[11][3] ) );
  XNOR2X1 U27 ( .A(\u_div/SumTmp[17][0] ), .B(\u_div/u_add_PartRem_1_11/n4 ), 
        .Y(\u_div/SumTmp[11][6] ) );
  NOR2X1 U28 ( .A(\u_div/u_add_PartRem_1_11/n4 ), .B(\u_div/SumTmp[17][0] ), 
        .Y(n14) );
  XOR2X1 U29 ( .A(\u_div/SumTmp[18][0] ), .B(n14), .Y(\u_div/SumTmp[11][7] )
         );
  NAND2BX1 U30 ( .AN(\u_div/SumTmp[18][0] ), .B(n14), .Y(
        \u_div/u_add_PartRem_1_11/n2 ) );
  CLKINVX1 U31 ( .A(\u_div/PartRem[11][3] ), .Y(\u_div/SumTmp[10][3] ) );
  XNOR2X1 U32 ( .A(\u_div/PartRem[11][6] ), .B(\u_div/u_add_PartRem_0_10/n5 ), 
        .Y(\u_div/SumTmp[10][6] ) );
  NOR2X1 U33 ( .A(\u_div/u_add_PartRem_0_10/n5 ), .B(\u_div/PartRem[11][6] ), 
        .Y(n15) );
  XOR2X1 U34 ( .A(\u_div/PartRem[11][7] ), .B(n15), .Y(\u_div/SumTmp[10][7] )
         );
  NAND2BX1 U35 ( .AN(\u_div/PartRem[11][7] ), .B(n15), .Y(
        \u_div/u_add_PartRem_0_10/n3 ) );
  CLKINVX1 U36 ( .A(\u_div/PartRem[10][3] ), .Y(\u_div/SumTmp[9][3] ) );
  XNOR2X1 U37 ( .A(\u_div/PartRem[10][6] ), .B(\u_div/u_add_PartRem_0_9/n5 ), 
        .Y(\u_div/SumTmp[9][6] ) );
  NOR2X1 U38 ( .A(\u_div/u_add_PartRem_0_9/n5 ), .B(\u_div/PartRem[10][6] ), 
        .Y(n16) );
  XOR2X1 U39 ( .A(\u_div/PartRem[10][7] ), .B(n16), .Y(\u_div/SumTmp[9][7] )
         );
  NAND2BX1 U40 ( .AN(\u_div/PartRem[10][7] ), .B(n16), .Y(
        \u_div/u_add_PartRem_0_9/n3 ) );
  CLKINVX1 U41 ( .A(\u_div/PartRem[9][3] ), .Y(\u_div/SumTmp[8][3] ) );
  XNOR2X1 U42 ( .A(\u_div/PartRem[9][6] ), .B(\u_div/u_add_PartRem_0_8/n5 ), 
        .Y(\u_div/SumTmp[8][6] ) );
  NOR2X1 U43 ( .A(\u_div/u_add_PartRem_0_8/n5 ), .B(\u_div/PartRem[9][6] ), 
        .Y(n17) );
  XOR2X1 U44 ( .A(\u_div/PartRem[9][7] ), .B(n17), .Y(\u_div/SumTmp[8][7] ) );
  NAND2BX1 U45 ( .AN(\u_div/PartRem[9][7] ), .B(n17), .Y(
        \u_div/u_add_PartRem_0_8/n3 ) );
  CLKINVX1 U46 ( .A(\u_div/PartRem[8][3] ), .Y(\u_div/SumTmp[7][3] ) );
  XNOR2X1 U47 ( .A(\u_div/PartRem[8][6] ), .B(\u_div/u_add_PartRem_0_7/n5 ), 
        .Y(\u_div/SumTmp[7][6] ) );
  NOR2X1 U48 ( .A(\u_div/u_add_PartRem_0_7/n5 ), .B(\u_div/PartRem[8][6] ), 
        .Y(n18) );
  XOR2X1 U49 ( .A(\u_div/PartRem[8][7] ), .B(n18), .Y(\u_div/SumTmp[7][7] ) );
  NAND2BX1 U50 ( .AN(\u_div/PartRem[8][7] ), .B(n18), .Y(
        \u_div/u_add_PartRem_0_7/n3 ) );
  CLKINVX1 U51 ( .A(\u_div/PartRem[7][3] ), .Y(\u_div/SumTmp[6][3] ) );
  XNOR2X1 U52 ( .A(\u_div/PartRem[7][6] ), .B(\u_div/u_add_PartRem_0_6/n5 ), 
        .Y(\u_div/SumTmp[6][6] ) );
  NOR2X1 U53 ( .A(\u_div/u_add_PartRem_0_6/n5 ), .B(\u_div/PartRem[7][6] ), 
        .Y(n19) );
  XOR2X1 U54 ( .A(\u_div/PartRem[7][7] ), .B(n19), .Y(\u_div/SumTmp[6][7] ) );
  NAND2BX1 U55 ( .AN(\u_div/PartRem[7][7] ), .B(n19), .Y(
        \u_div/u_add_PartRem_0_6/n3 ) );
  CLKINVX1 U56 ( .A(\u_div/PartRem[6][3] ), .Y(\u_div/SumTmp[5][3] ) );
  XNOR2X1 U57 ( .A(\u_div/PartRem[6][6] ), .B(\u_div/u_add_PartRem_0_5/n5 ), 
        .Y(\u_div/SumTmp[5][6] ) );
  NOR2X1 U58 ( .A(\u_div/u_add_PartRem_0_5/n5 ), .B(\u_div/PartRem[6][6] ), 
        .Y(n20) );
  XOR2X1 U59 ( .A(\u_div/PartRem[6][7] ), .B(n20), .Y(\u_div/SumTmp[5][7] ) );
  NAND2BX1 U60 ( .AN(\u_div/PartRem[6][7] ), .B(n20), .Y(
        \u_div/u_add_PartRem_0_5/n3 ) );
  CLKINVX1 U61 ( .A(\u_div/PartRem[5][3] ), .Y(\u_div/SumTmp[4][3] ) );
  XNOR2X1 U62 ( .A(\u_div/PartRem[5][6] ), .B(\u_div/u_add_PartRem_0_4/n5 ), 
        .Y(\u_div/SumTmp[4][6] ) );
  NOR2X1 U63 ( .A(\u_div/u_add_PartRem_0_4/n5 ), .B(\u_div/PartRem[5][6] ), 
        .Y(n21) );
  XOR2X1 U64 ( .A(\u_div/PartRem[5][7] ), .B(n21), .Y(\u_div/SumTmp[4][7] ) );
  NAND2BX1 U65 ( .AN(\u_div/PartRem[5][7] ), .B(n21), .Y(
        \u_div/u_add_PartRem_0_4/n3 ) );
  CLKINVX1 U66 ( .A(\u_div/PartRem[4][3] ), .Y(\u_div/SumTmp[3][3] ) );
  XNOR2X1 U67 ( .A(\u_div/PartRem[4][6] ), .B(\u_div/u_add_PartRem_0_3/n5 ), 
        .Y(\u_div/SumTmp[3][6] ) );
  NOR2X1 U68 ( .A(\u_div/u_add_PartRem_0_3/n5 ), .B(\u_div/PartRem[4][6] ), 
        .Y(n22) );
  XOR2X1 U69 ( .A(\u_div/PartRem[4][7] ), .B(n22), .Y(\u_div/SumTmp[3][7] ) );
  NAND2BX1 U70 ( .AN(\u_div/PartRem[4][7] ), .B(n22), .Y(
        \u_div/u_add_PartRem_0_3/n3 ) );
  CLKINVX1 U71 ( .A(\u_div/PartRem[3][3] ), .Y(\u_div/SumTmp[2][3] ) );
  XNOR2X1 U72 ( .A(\u_div/PartRem[3][6] ), .B(\u_div/u_add_PartRem_0_2/n5 ), 
        .Y(\u_div/SumTmp[2][6] ) );
  NOR2X1 U73 ( .A(\u_div/u_add_PartRem_0_2/n5 ), .B(\u_div/PartRem[3][6] ), 
        .Y(n23) );
  XOR2X1 U74 ( .A(\u_div/PartRem[3][7] ), .B(n23), .Y(\u_div/SumTmp[2][7] ) );
  NAND2BX1 U75 ( .AN(\u_div/PartRem[3][7] ), .B(n23), .Y(
        \u_div/u_add_PartRem_0_2/n3 ) );
  CLKINVX1 U76 ( .A(\u_div/PartRem[2][3] ), .Y(\u_div/SumTmp[1][3] ) );
  XNOR2X1 U77 ( .A(\u_div/PartRem[2][6] ), .B(\u_div/u_add_PartRem_0_1/n5 ), 
        .Y(\u_div/SumTmp[1][6] ) );
  NOR2X1 U78 ( .A(\u_div/u_add_PartRem_0_1/n5 ), .B(\u_div/PartRem[2][6] ), 
        .Y(n24) );
  XOR2X1 U79 ( .A(\u_div/PartRem[2][7] ), .B(n24), .Y(\u_div/SumTmp[1][7] ) );
  NAND2BX1 U80 ( .AN(\u_div/PartRem[2][7] ), .B(n24), .Y(
        \u_div/u_add_PartRem_0_1/n3 ) );
  OAI31XL U81 ( .A0(n25), .A1(\u_div/PartRem[1][7] ), .A2(
        \u_div/PartRem[1][6] ), .B0(\u_div/PartRem[1][8] ), .Y(n26) );
  NAND2BX1 U82 ( .AN(\u_div/PartRem[1][9] ), .B(n26), .Y(quotient[0]) );
endmodule


module CONT_DW_div_uns_12 ( a, b, quotient, remainder, divide_by_0 );
  input [31:0] a;
  input [2:0] b;
  output [31:0] quotient;
  output [2:0] remainder;
  output divide_by_0;
  wire   n87, \u_div/SumTmp[0][0] , \u_div/SumTmp[1][0] , \u_div/SumTmp[2][0] ,
         \u_div/SumTmp[3][0] , \u_div/SumTmp[4][0] , \u_div/SumTmp[5][0] ,
         \u_div/SumTmp[6][0] , \u_div/SumTmp[7][0] , \u_div/SumTmp[8][0] ,
         \u_div/SumTmp[9][0] , \u_div/SumTmp[10][0] , \u_div/SumTmp[11][0] ,
         \u_div/SumTmp[12][0] , \u_div/SumTmp[13][0] , \u_div/SumTmp[14][0] ,
         \u_div/SumTmp[15][0] , \u_div/SumTmp[16][0] , \u_div/SumTmp[17][0] ,
         \u_div/SumTmp[18][0] , \u_div/SumTmp[19][0] , n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86;
  assign \u_div/SumTmp[0][0]  = a[0];
  assign \u_div/SumTmp[1][0]  = a[1];
  assign \u_div/SumTmp[2][0]  = a[2];
  assign \u_div/SumTmp[3][0]  = a[3];
  assign \u_div/SumTmp[4][0]  = a[4];
  assign \u_div/SumTmp[5][0]  = a[5];
  assign \u_div/SumTmp[6][0]  = a[6];
  assign \u_div/SumTmp[7][0]  = a[7];
  assign \u_div/SumTmp[8][0]  = a[8];
  assign \u_div/SumTmp[9][0]  = a[9];
  assign \u_div/SumTmp[10][0]  = a[10];
  assign \u_div/SumTmp[11][0]  = a[11];
  assign \u_div/SumTmp[12][0]  = a[12];
  assign \u_div/SumTmp[13][0]  = a[13];
  assign \u_div/SumTmp[14][0]  = a[14];
  assign \u_div/SumTmp[15][0]  = a[15];
  assign \u_div/SumTmp[16][0]  = a[16];
  assign \u_div/SumTmp[17][0]  = a[17];
  assign \u_div/SumTmp[18][0]  = a[18];
  assign \u_div/SumTmp[19][0]  = a[19];

  MX2X1 \u_div/u_mx_PartRem_0_0_0  ( .A(\u_div/SumTmp[0][0] ), .B(
        \u_div/SumTmp[0][0] ), .S0(n1), .Y(remainder[0]) );
  OA21XL U1 ( .A0(n85), .A1(n84), .B0(n82), .Y(n87) );
  OA21X2 U2 ( .A0(n18), .A1(n19), .B0(n17), .Y(n21) );
  MXI2X1 U3 ( .A(n16), .B(n15), .S0(n14), .Y(n17) );
  OA21X2 U4 ( .A0(n33), .A1(n34), .B0(n32), .Y(n36) );
  MXI2X1 U5 ( .A(n31), .B(n30), .S0(n29), .Y(n32) );
  OA21X2 U6 ( .A0(n48), .A1(n49), .B0(n47), .Y(n51) );
  MXI2X1 U7 ( .A(n46), .B(n45), .S0(n44), .Y(n47) );
  OA21X2 U8 ( .A0(n63), .A1(n64), .B0(n62), .Y(n66) );
  MXI2X1 U9 ( .A(n61), .B(n60), .S0(n59), .Y(n62) );
  OA21X2 U10 ( .A0(n78), .A1(n79), .B0(n77), .Y(n81) );
  MXI2X1 U11 ( .A(n76), .B(n75), .S0(n74), .Y(n77) );
  OA21X2 U12 ( .A0(n13), .A1(n14), .B0(n12), .Y(n16) );
  MXI2X1 U13 ( .A(n11), .B(n10), .S0(n9), .Y(n12) );
  OA21X2 U14 ( .A0(n28), .A1(n29), .B0(n27), .Y(n31) );
  MXI2X1 U15 ( .A(n26), .B(n25), .S0(n24), .Y(n27) );
  OA21X2 U16 ( .A0(n43), .A1(n44), .B0(n42), .Y(n46) );
  MXI2X1 U17 ( .A(n41), .B(n40), .S0(n39), .Y(n42) );
  OA21X2 U18 ( .A0(n58), .A1(n59), .B0(n57), .Y(n61) );
  MXI2X1 U19 ( .A(n56), .B(n55), .S0(n54), .Y(n57) );
  OA21X2 U20 ( .A0(n73), .A1(n74), .B0(n72), .Y(n76) );
  MXI2X1 U21 ( .A(n71), .B(n70), .S0(n69), .Y(n72) );
  OA21X2 U22 ( .A0(n8), .A1(n9), .B0(n7), .Y(n11) );
  OA21X2 U23 ( .A0(n23), .A1(n24), .B0(n22), .Y(n26) );
  OA21X2 U24 ( .A0(n38), .A1(n39), .B0(n37), .Y(n41) );
  OA21X2 U25 ( .A0(n53), .A1(n54), .B0(n52), .Y(n56) );
  OA21X2 U26 ( .A0(n68), .A1(n69), .B0(n67), .Y(n71) );
  CLKINVX1 U27 ( .A(n87), .Y(n1) );
  XNOR2X2 U28 ( .A(n85), .B(n1), .Y(remainder[1]) );
  MXI2X2 U29 ( .A(n84), .B(n83), .S0(n1), .Y(remainder[2]) );
  MXI2XL U30 ( .A(n81), .B(n80), .S0(n79), .Y(n82) );
  NOR2XL U31 ( .A(n81), .B(n78), .Y(n80) );
  NOR2XL U32 ( .A(n76), .B(n73), .Y(n75) );
  NOR2XL U33 ( .A(n71), .B(n68), .Y(n70) );
  MXI2XL U34 ( .A(n66), .B(n65), .S0(n64), .Y(n67) );
  NOR2XL U35 ( .A(n66), .B(n63), .Y(n65) );
  NOR2XL U36 ( .A(n61), .B(n58), .Y(n60) );
  NOR2XL U37 ( .A(n56), .B(n53), .Y(n55) );
  MXI2XL U38 ( .A(n51), .B(n50), .S0(n49), .Y(n52) );
  NOR2XL U39 ( .A(n51), .B(n48), .Y(n50) );
  NOR2XL U40 ( .A(n46), .B(n43), .Y(n45) );
  NOR2XL U41 ( .A(n41), .B(n38), .Y(n40) );
  MXI2XL U42 ( .A(n36), .B(n35), .S0(n34), .Y(n37) );
  NOR2XL U43 ( .A(n36), .B(n33), .Y(n35) );
  NOR2XL U44 ( .A(n31), .B(n28), .Y(n30) );
  NOR2XL U45 ( .A(n26), .B(n23), .Y(n25) );
  MXI2XL U46 ( .A(n21), .B(n20), .S0(n19), .Y(n22) );
  NOR2XL U47 ( .A(n21), .B(n18), .Y(n20) );
  NOR2XL U48 ( .A(n16), .B(n13), .Y(n15) );
  NOR2XL U49 ( .A(n11), .B(n8), .Y(n10) );
  CLKINVX1 U50 ( .A(\u_div/SumTmp[18][0] ), .Y(n86) );
  CLKINVX1 U51 ( .A(\u_div/SumTmp[1][0] ), .Y(n85) );
  CLKINVX1 U52 ( .A(\u_div/SumTmp[2][0] ), .Y(n78) );
  CLKINVX1 U53 ( .A(\u_div/SumTmp[3][0] ), .Y(n73) );
  CLKINVX1 U54 ( .A(\u_div/SumTmp[4][0] ), .Y(n68) );
  CLKINVX1 U55 ( .A(\u_div/SumTmp[5][0] ), .Y(n63) );
  CLKINVX1 U56 ( .A(\u_div/SumTmp[6][0] ), .Y(n58) );
  CLKINVX1 U57 ( .A(\u_div/SumTmp[7][0] ), .Y(n53) );
  CLKINVX1 U58 ( .A(\u_div/SumTmp[8][0] ), .Y(n48) );
  CLKINVX1 U59 ( .A(\u_div/SumTmp[9][0] ), .Y(n43) );
  CLKINVX1 U60 ( .A(\u_div/SumTmp[10][0] ), .Y(n38) );
  CLKINVX1 U61 ( .A(\u_div/SumTmp[11][0] ), .Y(n33) );
  CLKINVX1 U62 ( .A(\u_div/SumTmp[12][0] ), .Y(n28) );
  CLKINVX1 U63 ( .A(\u_div/SumTmp[13][0] ), .Y(n23) );
  CLKINVX1 U64 ( .A(\u_div/SumTmp[14][0] ), .Y(n18) );
  CLKINVX1 U65 ( .A(\u_div/SumTmp[15][0] ), .Y(n13) );
  CLKINVX1 U66 ( .A(\u_div/SumTmp[16][0] ), .Y(n8) );
  CLKINVX1 U67 ( .A(\u_div/SumTmp[17][0] ), .Y(n3) );
  NAND2X1 U68 ( .A(\u_div/SumTmp[18][0] ), .B(\u_div/SumTmp[19][0] ), .Y(n2)
         );
  MXI2X1 U69 ( .A(n86), .B(\u_div/SumTmp[18][0] ), .S0(n2), .Y(n4) );
  AOI2BB2X1 U70 ( .B0(n2), .B1(\u_div/SumTmp[19][0] ), .A0N(n4), .A1N(n3), .Y(
        n6) );
  XNOR2X1 U71 ( .A(n3), .B(n6), .Y(n9) );
  NOR2X1 U72 ( .A(n6), .B(n3), .Y(n5) );
  MXI2X1 U73 ( .A(n6), .B(n5), .S0(n4), .Y(n7) );
  XNOR2X1 U74 ( .A(n8), .B(n11), .Y(n14) );
  XNOR2X1 U75 ( .A(n13), .B(n16), .Y(n19) );
  XNOR2X1 U76 ( .A(n18), .B(n21), .Y(n24) );
  XNOR2X1 U77 ( .A(n23), .B(n26), .Y(n29) );
  XNOR2X1 U78 ( .A(n28), .B(n31), .Y(n34) );
  XNOR2X1 U79 ( .A(n33), .B(n36), .Y(n39) );
  XNOR2X1 U80 ( .A(n38), .B(n41), .Y(n44) );
  XNOR2X1 U81 ( .A(n43), .B(n46), .Y(n49) );
  XNOR2X1 U82 ( .A(n48), .B(n51), .Y(n54) );
  XNOR2X1 U83 ( .A(n53), .B(n56), .Y(n59) );
  XNOR2X1 U84 ( .A(n58), .B(n61), .Y(n64) );
  XNOR2X1 U85 ( .A(n63), .B(n66), .Y(n69) );
  XNOR2X1 U86 ( .A(n68), .B(n71), .Y(n74) );
  XNOR2X1 U87 ( .A(n73), .B(n76), .Y(n79) );
  XNOR2X1 U88 ( .A(n78), .B(n81), .Y(n84) );
  NAND2X1 U89 ( .A(\u_div/SumTmp[1][0] ), .B(n84), .Y(n83) );
endmodule


module CONT_DW_div_uns_13 ( a, b, quotient, remainder, divide_by_0 );
  input [31:0] a;
  input [3:0] b;
  output [31:0] quotient;
  output [3:0] remainder;
  output divide_by_0;
  wire   n130, \u_div/SumTmp[0][0] , \u_div/SumTmp[1][0] ,
         \u_div/SumTmp[2][0] , \u_div/SumTmp[3][0] , \u_div/SumTmp[4][0] ,
         \u_div/SumTmp[5][0] , \u_div/SumTmp[6][0] , \u_div/SumTmp[7][0] ,
         \u_div/SumTmp[8][0] , \u_div/SumTmp[9][0] , \u_div/SumTmp[10][0] ,
         \u_div/SumTmp[11][0] , \u_div/SumTmp[12][0] , \u_div/SumTmp[13][0] ,
         \u_div/SumTmp[14][0] , \u_div/SumTmp[15][0] , \u_div/SumTmp[16][0] ,
         \u_div/SumTmp[16][2] , \u_div/SumTmp[17][0] , \u_div/SumTmp[18][0] ,
         \u_div/SumTmp[19][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129;
  assign \u_div/SumTmp[0][0]  = a[0];
  assign \u_div/SumTmp[1][0]  = a[1];
  assign \u_div/SumTmp[2][0]  = a[2];
  assign \u_div/SumTmp[3][0]  = a[3];
  assign \u_div/SumTmp[4][0]  = a[4];
  assign \u_div/SumTmp[5][0]  = a[5];
  assign \u_div/SumTmp[6][0]  = a[6];
  assign \u_div/SumTmp[7][0]  = a[7];
  assign \u_div/SumTmp[8][0]  = a[8];
  assign \u_div/SumTmp[9][0]  = a[9];
  assign \u_div/SumTmp[10][0]  = a[10];
  assign \u_div/SumTmp[11][0]  = a[11];
  assign \u_div/SumTmp[12][0]  = a[12];
  assign \u_div/SumTmp[13][0]  = a[13];
  assign \u_div/SumTmp[14][0]  = a[14];
  assign \u_div/SumTmp[15][0]  = a[15];
  assign \u_div/SumTmp[16][0]  = a[16];
  assign \u_div/SumTmp[17][0]  = a[17];
  assign \u_div/SumTmp[18][0]  = a[18];
  assign \u_div/SumTmp[19][0]  = a[19];

  MX2XL \u_div/u_mx_PartRem_0_0_0  ( .A(\u_div/SumTmp[0][0] ), .B(
        \u_div/SumTmp[0][0] ), .S0(n130), .Y(remainder[0]) );
  OA21X2 U1 ( .A0(n100), .A1(n101), .B0(n97), .Y(n102) );
  AOI2BB2X2 U2 ( .B0(n1), .B1(\u_div/SumTmp[19][0] ), .A0N(n4), .A1N(n5), .Y(
        n6) );
  OA21X2 U3 ( .A0(n76), .A1(n77), .B0(n73), .Y(n78) );
  OA21X2 U4 ( .A0(n52), .A1(n53), .B0(n49), .Y(n54) );
  OA21X2 U5 ( .A0(n28), .A1(n29), .B0(n25), .Y(n30) );
  OA21X2 U6 ( .A0(n108), .A1(n109), .B0(n105), .Y(n110) );
  OA21X2 U7 ( .A0(n12), .A1(n13), .B0(n9), .Y(n14) );
  OA21X2 U8 ( .A0(n84), .A1(n85), .B0(n81), .Y(n86) );
  OA21X2 U9 ( .A0(n60), .A1(n61), .B0(n57), .Y(n62) );
  OA21X2 U10 ( .A0(n36), .A1(n37), .B0(n33), .Y(n38) );
  MXI2X2 U11 ( .A(n115), .B(n114), .S0(n118), .Y(n124) );
  OA21X2 U12 ( .A0(n92), .A1(n93), .B0(n89), .Y(n94) );
  OA21X2 U13 ( .A0(n68), .A1(n69), .B0(n65), .Y(n70) );
  OA21X2 U14 ( .A0(n44), .A1(n45), .B0(n41), .Y(n46) );
  OA21X2 U15 ( .A0(n20), .A1(n21), .B0(n17), .Y(n22) );
  OAI21X2 U16 ( .A0(n124), .A1(n122), .B0(n121), .Y(n130) );
  OA21X2 U17 ( .A0(n116), .A1(n117), .B0(n113), .Y(n118) );
  MXI2XL U18 ( .A(n120), .B(n119), .S0(n118), .Y(n121) );
  MXI2XL U19 ( .A(n104), .B(n103), .S0(n102), .Y(n105) );
  MXI2XL U20 ( .A(n64), .B(n63), .S0(n62), .Y(n65) );
  MXI2XL U21 ( .A(n112), .B(n111), .S0(n110), .Y(n113) );
  MXI2XL U22 ( .A(n124), .B(n123), .S0(n130), .Y(remainder[3]) );
  XNOR2XL U23 ( .A(n122), .B(n124), .Y(n123) );
  MXI2XL U24 ( .A(n127), .B(n126), .S0(n130), .Y(remainder[2]) );
  XNOR2XL U25 ( .A(n125), .B(n130), .Y(remainder[1]) );
  MXI2XL U26 ( .A(n96), .B(n95), .S0(n94), .Y(n97) );
  MXI2XL U27 ( .A(n8), .B(n7), .S0(n6), .Y(n9) );
  MXI2XL U28 ( .A(n16), .B(n15), .S0(n14), .Y(n17) );
  MXI2XL U29 ( .A(n24), .B(n23), .S0(n22), .Y(n25) );
  MXI2XL U30 ( .A(n32), .B(n31), .S0(n30), .Y(n33) );
  MXI2XL U31 ( .A(n40), .B(n39), .S0(n38), .Y(n41) );
  MXI2XL U32 ( .A(n48), .B(n47), .S0(n46), .Y(n49) );
  MXI2XL U33 ( .A(n56), .B(n55), .S0(n54), .Y(n57) );
  MXI2XL U34 ( .A(n72), .B(n71), .S0(n70), .Y(n73) );
  MXI2XL U35 ( .A(n80), .B(n79), .S0(n78), .Y(n81) );
  MXI2XL U36 ( .A(n88), .B(n87), .S0(n86), .Y(n89) );
  CLKINVX1 U37 ( .A(\u_div/SumTmp[17][0] ), .Y(n128) );
  NAND2X1 U38 ( .A(n129), .B(\u_div/SumTmp[19][0] ), .Y(n1) );
  CLKMX2X2 U39 ( .A(n128), .B(\u_div/SumTmp[17][0] ), .S0(n1), .Y(n2) );
  XOR2X1 U40 ( .A(\u_div/SumTmp[16][0] ), .B(n2), .Y(n3) );
  MXI2X1 U41 ( .A(\u_div/SumTmp[16][2] ), .B(\u_div/SumTmp[18][0] ), .S0(n1), 
        .Y(n4) );
  NAND2X1 U42 ( .A(\u_div/SumTmp[16][0] ), .B(n2), .Y(n5) );
  MXI2X1 U43 ( .A(n3), .B(n2), .S0(n6), .Y(n12) );
  XNOR2X1 U44 ( .A(\u_div/SumTmp[16][0] ), .B(n6), .Y(n10) );
  NAND2X1 U45 ( .A(\u_div/SumTmp[15][0] ), .B(n10), .Y(n13) );
  CLKINVX1 U46 ( .A(n4), .Y(n7) );
  XNOR2X1 U47 ( .A(n5), .B(n7), .Y(n8) );
  XNOR2X1 U48 ( .A(\u_div/SumTmp[15][0] ), .B(n14), .Y(n18) );
  XOR2X1 U49 ( .A(n18), .B(\u_div/SumTmp[14][0] ), .Y(n19) );
  XOR2X1 U50 ( .A(n10), .B(\u_div/SumTmp[15][0] ), .Y(n11) );
  MXI2X1 U51 ( .A(n11), .B(n10), .S0(n14), .Y(n20) );
  NAND2X1 U52 ( .A(\u_div/SumTmp[14][0] ), .B(n18), .Y(n21) );
  CLKINVX1 U53 ( .A(n12), .Y(n15) );
  XNOR2X1 U54 ( .A(n13), .B(n15), .Y(n16) );
  MXI2X1 U55 ( .A(n19), .B(n18), .S0(n22), .Y(n28) );
  XNOR2X1 U56 ( .A(\u_div/SumTmp[14][0] ), .B(n22), .Y(n26) );
  NAND2X1 U57 ( .A(\u_div/SumTmp[13][0] ), .B(n26), .Y(n29) );
  CLKINVX1 U58 ( .A(n20), .Y(n23) );
  XNOR2X1 U59 ( .A(n21), .B(n23), .Y(n24) );
  XNOR2X1 U60 ( .A(\u_div/SumTmp[13][0] ), .B(n30), .Y(n34) );
  XOR2X1 U61 ( .A(n34), .B(\u_div/SumTmp[12][0] ), .Y(n35) );
  XOR2X1 U62 ( .A(n26), .B(\u_div/SumTmp[13][0] ), .Y(n27) );
  MXI2X1 U63 ( .A(n27), .B(n26), .S0(n30), .Y(n36) );
  NAND2X1 U64 ( .A(\u_div/SumTmp[12][0] ), .B(n34), .Y(n37) );
  CLKINVX1 U65 ( .A(n28), .Y(n31) );
  XNOR2X1 U66 ( .A(n29), .B(n31), .Y(n32) );
  MXI2X1 U67 ( .A(n35), .B(n34), .S0(n38), .Y(n44) );
  XNOR2X1 U68 ( .A(\u_div/SumTmp[12][0] ), .B(n38), .Y(n42) );
  NAND2X1 U69 ( .A(\u_div/SumTmp[11][0] ), .B(n42), .Y(n45) );
  CLKINVX1 U70 ( .A(n36), .Y(n39) );
  XNOR2X1 U71 ( .A(n37), .B(n39), .Y(n40) );
  XNOR2X1 U72 ( .A(\u_div/SumTmp[11][0] ), .B(n46), .Y(n50) );
  XOR2X1 U73 ( .A(n50), .B(\u_div/SumTmp[10][0] ), .Y(n51) );
  XOR2X1 U74 ( .A(n42), .B(\u_div/SumTmp[11][0] ), .Y(n43) );
  MXI2X1 U75 ( .A(n43), .B(n42), .S0(n46), .Y(n52) );
  NAND2X1 U76 ( .A(\u_div/SumTmp[10][0] ), .B(n50), .Y(n53) );
  CLKINVX1 U77 ( .A(n44), .Y(n47) );
  XNOR2X1 U78 ( .A(n45), .B(n47), .Y(n48) );
  MXI2X1 U79 ( .A(n51), .B(n50), .S0(n54), .Y(n60) );
  XNOR2X1 U80 ( .A(\u_div/SumTmp[10][0] ), .B(n54), .Y(n58) );
  NAND2X1 U81 ( .A(\u_div/SumTmp[9][0] ), .B(n58), .Y(n61) );
  CLKINVX1 U82 ( .A(n52), .Y(n55) );
  XNOR2X1 U83 ( .A(n53), .B(n55), .Y(n56) );
  XNOR2X1 U84 ( .A(\u_div/SumTmp[9][0] ), .B(n62), .Y(n66) );
  XOR2X1 U85 ( .A(n66), .B(\u_div/SumTmp[8][0] ), .Y(n67) );
  XOR2X1 U86 ( .A(n58), .B(\u_div/SumTmp[9][0] ), .Y(n59) );
  MXI2X1 U87 ( .A(n59), .B(n58), .S0(n62), .Y(n68) );
  NAND2X1 U88 ( .A(\u_div/SumTmp[8][0] ), .B(n66), .Y(n69) );
  CLKINVX1 U89 ( .A(n60), .Y(n63) );
  XNOR2X1 U90 ( .A(n61), .B(n63), .Y(n64) );
  MXI2X1 U91 ( .A(n67), .B(n66), .S0(n70), .Y(n76) );
  XNOR2X1 U92 ( .A(\u_div/SumTmp[8][0] ), .B(n70), .Y(n74) );
  NAND2X1 U93 ( .A(\u_div/SumTmp[7][0] ), .B(n74), .Y(n77) );
  CLKINVX1 U94 ( .A(n68), .Y(n71) );
  XNOR2X1 U95 ( .A(n69), .B(n71), .Y(n72) );
  XNOR2X1 U96 ( .A(\u_div/SumTmp[7][0] ), .B(n78), .Y(n82) );
  XOR2X1 U97 ( .A(n82), .B(\u_div/SumTmp[6][0] ), .Y(n83) );
  XOR2X1 U98 ( .A(n74), .B(\u_div/SumTmp[7][0] ), .Y(n75) );
  MXI2X1 U99 ( .A(n75), .B(n74), .S0(n78), .Y(n84) );
  NAND2X1 U100 ( .A(\u_div/SumTmp[6][0] ), .B(n82), .Y(n85) );
  CLKINVX1 U101 ( .A(n76), .Y(n79) );
  XNOR2X1 U102 ( .A(n77), .B(n79), .Y(n80) );
  MXI2X1 U103 ( .A(n83), .B(n82), .S0(n86), .Y(n92) );
  XNOR2X1 U104 ( .A(\u_div/SumTmp[6][0] ), .B(n86), .Y(n90) );
  NAND2X1 U105 ( .A(\u_div/SumTmp[5][0] ), .B(n90), .Y(n93) );
  CLKINVX1 U106 ( .A(n84), .Y(n87) );
  XNOR2X1 U107 ( .A(n85), .B(n87), .Y(n88) );
  XNOR2X1 U108 ( .A(\u_div/SumTmp[5][0] ), .B(n94), .Y(n98) );
  XOR2X1 U109 ( .A(n98), .B(\u_div/SumTmp[4][0] ), .Y(n99) );
  XOR2X1 U110 ( .A(n90), .B(\u_div/SumTmp[5][0] ), .Y(n91) );
  MXI2X1 U111 ( .A(n91), .B(n90), .S0(n94), .Y(n100) );
  NAND2X1 U112 ( .A(\u_div/SumTmp[4][0] ), .B(n98), .Y(n101) );
  CLKINVX1 U113 ( .A(n92), .Y(n95) );
  XNOR2X1 U114 ( .A(n93), .B(n95), .Y(n96) );
  MXI2X1 U115 ( .A(n99), .B(n98), .S0(n102), .Y(n108) );
  XNOR2X1 U116 ( .A(\u_div/SumTmp[4][0] ), .B(n102), .Y(n106) );
  NAND2X1 U117 ( .A(\u_div/SumTmp[3][0] ), .B(n106), .Y(n109) );
  CLKINVX1 U118 ( .A(n100), .Y(n103) );
  XNOR2X1 U119 ( .A(n101), .B(n103), .Y(n104) );
  XNOR2X1 U120 ( .A(\u_div/SumTmp[3][0] ), .B(n110), .Y(n114) );
  XOR2X1 U121 ( .A(n114), .B(\u_div/SumTmp[2][0] ), .Y(n115) );
  XOR2X1 U122 ( .A(n106), .B(\u_div/SumTmp[3][0] ), .Y(n107) );
  MXI2X1 U123 ( .A(n107), .B(n106), .S0(n110), .Y(n116) );
  NAND2X1 U124 ( .A(\u_div/SumTmp[2][0] ), .B(n114), .Y(n117) );
  CLKINVX1 U125 ( .A(n108), .Y(n111) );
  XNOR2X1 U126 ( .A(n109), .B(n111), .Y(n112) );
  XOR2X1 U127 ( .A(\u_div/SumTmp[2][0] ), .B(n118), .Y(n127) );
  NAND2BX1 U128 ( .AN(n127), .B(\u_div/SumTmp[1][0] ), .Y(n122) );
  CLKINVX1 U129 ( .A(n116), .Y(n119) );
  XNOR2X1 U130 ( .A(n117), .B(n119), .Y(n120) );
  CLKINVX1 U131 ( .A(\u_div/SumTmp[1][0] ), .Y(n125) );
  XNOR2X1 U132 ( .A(n125), .B(n127), .Y(n126) );
  NOR2BX1 U133 ( .AN(\u_div/SumTmp[18][0] ), .B(n128), .Y(n129) );
  XOR2X1 U134 ( .A(\u_div/SumTmp[18][0] ), .B(\u_div/SumTmp[17][0] ), .Y(
        \u_div/SumTmp[16][2] ) );
endmodule


module CONT_DW_div_uns_14 ( a, b, quotient, remainder, divide_by_0 );
  input [20:0] a;
  input [2:0] b;
  output [20:0] quotient;
  output [2:0] remainder;
  output divide_by_0;
  wire   n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, \u_div/SumTmp[0][1] , \u_div/SumTmp[0][2] ,
         \u_div/SumTmp[1][1] , \u_div/SumTmp[1][2] , \u_div/SumTmp[2][1] ,
         \u_div/SumTmp[2][2] , \u_div/SumTmp[3][1] , \u_div/SumTmp[3][2] ,
         \u_div/SumTmp[4][1] , \u_div/SumTmp[4][2] , \u_div/SumTmp[5][1] ,
         \u_div/SumTmp[5][2] , \u_div/SumTmp[6][1] , \u_div/SumTmp[6][2] ,
         \u_div/SumTmp[7][1] , \u_div/SumTmp[7][2] , \u_div/SumTmp[8][1] ,
         \u_div/SumTmp[8][2] , \u_div/SumTmp[9][1] , \u_div/SumTmp[9][2] ,
         \u_div/SumTmp[10][1] , \u_div/SumTmp[10][2] , \u_div/SumTmp[11][1] ,
         \u_div/SumTmp[11][2] , \u_div/SumTmp[12][1] , \u_div/SumTmp[12][2] ,
         \u_div/SumTmp[13][1] , \u_div/SumTmp[13][2] , \u_div/SumTmp[14][1] ,
         \u_div/SumTmp[14][2] , \u_div/SumTmp[15][1] , \u_div/SumTmp[15][2] ,
         \u_div/SumTmp[16][1] , \u_div/SumTmp[16][2] , \u_div/SumTmp[17][1] ,
         \u_div/SumTmp[17][2] , \u_div/SumTmp[18][1] , \u_div/SumTmp[18][2] ,
         \u_div/CryTmp[0][1] , \u_div/CryTmp[1][1] , \u_div/CryTmp[2][1] ,
         \u_div/CryTmp[3][1] , \u_div/CryTmp[4][1] , \u_div/CryTmp[5][1] ,
         \u_div/CryTmp[6][1] , \u_div/CryTmp[7][1] , \u_div/CryTmp[8][1] ,
         \u_div/CryTmp[9][1] , \u_div/CryTmp[10][1] , \u_div/CryTmp[11][1] ,
         \u_div/CryTmp[12][1] , \u_div/CryTmp[13][1] , \u_div/CryTmp[14][1] ,
         \u_div/CryTmp[15][1] , \u_div/CryTmp[16][1] , \u_div/CryTmp[17][1] ,
         \u_div/CryTmp[18][1] , \u_div/CryTmp[19][1] , \u_div/PartRem[1][1] ,
         \u_div/PartRem[1][2] , \u_div/PartRem[2][1] , \u_div/PartRem[2][2] ,
         \u_div/PartRem[3][1] , \u_div/PartRem[3][2] , \u_div/PartRem[4][1] ,
         \u_div/PartRem[4][2] , \u_div/PartRem[5][1] , \u_div/PartRem[5][2] ,
         \u_div/PartRem[6][1] , \u_div/PartRem[6][2] , \u_div/PartRem[7][1] ,
         \u_div/PartRem[7][2] , \u_div/PartRem[8][1] , \u_div/PartRem[8][2] ,
         \u_div/PartRem[9][1] , \u_div/PartRem[9][2] , \u_div/PartRem[10][1] ,
         \u_div/PartRem[10][2] , \u_div/PartRem[11][1] ,
         \u_div/PartRem[11][2] , \u_div/PartRem[12][1] ,
         \u_div/PartRem[12][2] , \u_div/PartRem[13][1] ,
         \u_div/PartRem[13][2] , \u_div/PartRem[14][1] ,
         \u_div/PartRem[14][2] , \u_div/PartRem[15][1] ,
         \u_div/PartRem[15][2] , \u_div/PartRem[16][1] ,
         \u_div/PartRem[16][2] , \u_div/PartRem[17][1] ,
         \u_div/PartRem[17][2] , \u_div/PartRem[18][1] ,
         \u_div/PartRem[18][2] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56;
  assign \u_div/CryTmp[0][1]  = a[0];
  assign \u_div/CryTmp[1][1]  = a[1];
  assign \u_div/CryTmp[2][1]  = a[2];
  assign \u_div/CryTmp[3][1]  = a[3];
  assign \u_div/CryTmp[4][1]  = a[4];
  assign \u_div/CryTmp[5][1]  = a[5];
  assign \u_div/CryTmp[6][1]  = a[6];
  assign \u_div/CryTmp[7][1]  = a[7];
  assign \u_div/CryTmp[8][1]  = a[8];
  assign \u_div/CryTmp[9][1]  = a[9];
  assign \u_div/CryTmp[10][1]  = a[10];
  assign \u_div/CryTmp[11][1]  = a[11];
  assign \u_div/CryTmp[12][1]  = a[12];
  assign \u_div/CryTmp[13][1]  = a[13];
  assign \u_div/CryTmp[14][1]  = a[14];
  assign \u_div/CryTmp[15][1]  = a[15];
  assign \u_div/CryTmp[16][1]  = a[16];
  assign \u_div/CryTmp[17][1]  = a[17];
  assign \u_div/CryTmp[18][1]  = a[18];
  assign \u_div/CryTmp[19][1]  = a[19];

  CLKMX2X2 \u_div/u_mx_PartRem_0_4_1  ( .A(\u_div/PartRem[5][1] ), .B(
        \u_div/SumTmp[4][1] ), .S0(n71), .Y(\u_div/PartRem[4][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_5_1  ( .A(\u_div/PartRem[6][1] ), .B(
        \u_div/SumTmp[5][1] ), .S0(n70), .Y(\u_div/PartRem[5][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_6_1  ( .A(\u_div/PartRem[7][1] ), .B(
        \u_div/SumTmp[6][1] ), .S0(n69), .Y(\u_div/PartRem[6][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_7_1  ( .A(\u_div/PartRem[8][1] ), .B(
        \u_div/SumTmp[7][1] ), .S0(n68), .Y(\u_div/PartRem[7][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_8_1  ( .A(\u_div/PartRem[9][1] ), .B(
        \u_div/SumTmp[8][1] ), .S0(n67), .Y(\u_div/PartRem[8][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_9_1  ( .A(\u_div/PartRem[10][1] ), .B(
        \u_div/SumTmp[9][1] ), .S0(n66), .Y(\u_div/PartRem[9][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_10_1  ( .A(\u_div/PartRem[11][1] ), .B(
        \u_div/SumTmp[10][1] ), .S0(n65), .Y(\u_div/PartRem[10][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_11_1  ( .A(\u_div/PartRem[12][1] ), .B(
        \u_div/SumTmp[11][1] ), .S0(n64), .Y(\u_div/PartRem[11][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_12_1  ( .A(\u_div/PartRem[13][1] ), .B(
        \u_div/SumTmp[12][1] ), .S0(n63), .Y(\u_div/PartRem[12][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_13_1  ( .A(\u_div/PartRem[14][1] ), .B(
        \u_div/SumTmp[13][1] ), .S0(n62), .Y(\u_div/PartRem[13][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_14_1  ( .A(\u_div/PartRem[15][1] ), .B(
        \u_div/SumTmp[14][1] ), .S0(n61), .Y(\u_div/PartRem[14][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_15_1  ( .A(\u_div/PartRem[16][1] ), .B(
        \u_div/SumTmp[15][1] ), .S0(n60), .Y(\u_div/PartRem[15][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_16_1  ( .A(\u_div/PartRem[17][1] ), .B(
        \u_div/SumTmp[16][1] ), .S0(n59), .Y(\u_div/PartRem[16][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_17_1  ( .A(\u_div/PartRem[18][1] ), .B(
        \u_div/SumTmp[17][1] ), .S0(n58), .Y(\u_div/PartRem[17][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_4_0  ( .A(\u_div/CryTmp[4][1] ), .B(n34), 
        .S0(n71), .Y(\u_div/PartRem[4][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_5_0  ( .A(\u_div/CryTmp[5][1] ), .B(n33), 
        .S0(n70), .Y(\u_div/PartRem[5][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_6_0  ( .A(\u_div/CryTmp[6][1] ), .B(n32), 
        .S0(n69), .Y(\u_div/PartRem[6][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_7_0  ( .A(\u_div/CryTmp[7][1] ), .B(n31), 
        .S0(n68), .Y(\u_div/PartRem[7][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_8_0  ( .A(\u_div/CryTmp[8][1] ), .B(n30), 
        .S0(n67), .Y(\u_div/PartRem[8][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_9_0  ( .A(\u_div/CryTmp[9][1] ), .B(n29), 
        .S0(n66), .Y(\u_div/PartRem[9][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_10_0  ( .A(\u_div/CryTmp[10][1] ), .B(n28), 
        .S0(n65), .Y(\u_div/PartRem[10][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_11_0  ( .A(\u_div/CryTmp[11][1] ), .B(n27), 
        .S0(n64), .Y(\u_div/PartRem[11][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_12_0  ( .A(\u_div/CryTmp[12][1] ), .B(n26), 
        .S0(n63), .Y(\u_div/PartRem[12][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_13_0  ( .A(\u_div/CryTmp[13][1] ), .B(n25), 
        .S0(n62), .Y(\u_div/PartRem[13][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_14_0  ( .A(\u_div/CryTmp[14][1] ), .B(n24), 
        .S0(n61), .Y(\u_div/PartRem[14][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_15_0  ( .A(\u_div/CryTmp[15][1] ), .B(n23), 
        .S0(n60), .Y(\u_div/PartRem[15][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_16_0  ( .A(\u_div/CryTmp[16][1] ), .B(n22), 
        .S0(n59), .Y(\u_div/PartRem[16][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_17_0  ( .A(\u_div/CryTmp[17][1] ), .B(n21), 
        .S0(n58), .Y(\u_div/PartRem[17][1] ) );
  MX2X1 \u_div/u_mx_PartRem_0_18_1  ( .A(\u_div/CryTmp[19][1] ), .B(
        \u_div/SumTmp[18][1] ), .S0(n57), .Y(\u_div/PartRem[18][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_18_0  ( .A(\u_div/CryTmp[18][1] ), .B(n20), .S0(
        n57), .Y(\u_div/PartRem[18][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_1_1  ( .A(\u_div/PartRem[2][1] ), .B(
        \u_div/SumTmp[1][1] ), .S0(n74), .Y(\u_div/PartRem[1][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_2_1  ( .A(\u_div/PartRem[3][1] ), .B(
        \u_div/SumTmp[2][1] ), .S0(n73), .Y(\u_div/PartRem[2][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_3_1  ( .A(\u_div/PartRem[4][1] ), .B(
        \u_div/SumTmp[3][1] ), .S0(n72), .Y(\u_div/PartRem[3][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_1_0  ( .A(\u_div/CryTmp[1][1] ), .B(n37), 
        .S0(n74), .Y(\u_div/PartRem[1][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_2_0  ( .A(\u_div/CryTmp[2][1] ), .B(n36), 
        .S0(n73), .Y(\u_div/PartRem[2][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_3_0  ( .A(\u_div/CryTmp[3][1] ), .B(n35), 
        .S0(n72), .Y(\u_div/PartRem[3][1] ) );
  MX2XL \u_div/u_mx_PartRem_0_0_0  ( .A(\u_div/CryTmp[0][1] ), .B(n19), .S0(
        n75), .Y(remainder[0]) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_0_2  ( .A(\u_div/PartRem[1][2] ), .B(
        \u_div/SumTmp[0][2] ), .S0(n75), .Y(remainder[2]) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_0_1  ( .A(\u_div/PartRem[1][1] ), .B(
        \u_div/SumTmp[0][1] ), .S0(n75), .Y(remainder[1]) );
  OR2XL U1 ( .A(\u_div/CryTmp[0][1] ), .B(\u_div/PartRem[1][1] ), .Y(n38) );
  XNOR2XL U2 ( .A(\u_div/PartRem[1][1] ), .B(\u_div/CryTmp[0][1] ), .Y(
        \u_div/SumTmp[0][1] ) );
  OAI2BB1X1 U3 ( .A0N(\u_div/PartRem[2][2] ), .A1N(n39), .B0(n1), .Y(n74) );
  MXI2X1 U4 ( .A(\u_div/PartRem[3][2] ), .B(\u_div/SumTmp[2][2] ), .S0(n73), 
        .Y(n1) );
  OAI2BB1X1 U5 ( .A0N(\u_div/PartRem[1][2] ), .A1N(n38), .B0(n2), .Y(n75) );
  MXI2X1 U6 ( .A(\u_div/PartRem[2][2] ), .B(\u_div/SumTmp[1][2] ), .S0(n74), 
        .Y(n2) );
  OAI2BB1X1 U7 ( .A0N(\u_div/PartRem[17][2] ), .A1N(n54), .B0(n3), .Y(n59) );
  MXI2X1 U8 ( .A(\u_div/PartRem[18][2] ), .B(\u_div/SumTmp[17][2] ), .S0(n58), 
        .Y(n3) );
  OAI2BB1X1 U9 ( .A0N(\u_div/PartRem[16][2] ), .A1N(n53), .B0(n4), .Y(n60) );
  MXI2X1 U10 ( .A(\u_div/PartRem[17][2] ), .B(\u_div/SumTmp[16][2] ), .S0(n59), 
        .Y(n4) );
  OAI2BB1X1 U11 ( .A0N(\u_div/PartRem[15][2] ), .A1N(n52), .B0(n5), .Y(n61) );
  MXI2X1 U12 ( .A(\u_div/PartRem[16][2] ), .B(\u_div/SumTmp[15][2] ), .S0(n60), 
        .Y(n5) );
  OAI2BB1X1 U13 ( .A0N(\u_div/PartRem[14][2] ), .A1N(n51), .B0(n6), .Y(n62) );
  MXI2X1 U14 ( .A(\u_div/PartRem[15][2] ), .B(\u_div/SumTmp[14][2] ), .S0(n61), 
        .Y(n6) );
  OAI2BB1X1 U15 ( .A0N(\u_div/PartRem[13][2] ), .A1N(n50), .B0(n7), .Y(n63) );
  MXI2X1 U16 ( .A(\u_div/PartRem[14][2] ), .B(\u_div/SumTmp[13][2] ), .S0(n62), 
        .Y(n7) );
  OAI2BB1X1 U17 ( .A0N(\u_div/PartRem[12][2] ), .A1N(n49), .B0(n8), .Y(n64) );
  MXI2X1 U18 ( .A(\u_div/PartRem[13][2] ), .B(\u_div/SumTmp[12][2] ), .S0(n63), 
        .Y(n8) );
  OAI2BB1X1 U19 ( .A0N(\u_div/PartRem[11][2] ), .A1N(n48), .B0(n9), .Y(n65) );
  MXI2X1 U20 ( .A(\u_div/PartRem[12][2] ), .B(\u_div/SumTmp[11][2] ), .S0(n64), 
        .Y(n9) );
  OAI2BB1X1 U21 ( .A0N(\u_div/PartRem[10][2] ), .A1N(n47), .B0(n10), .Y(n66)
         );
  MXI2X1 U22 ( .A(\u_div/PartRem[11][2] ), .B(\u_div/SumTmp[10][2] ), .S0(n65), 
        .Y(n10) );
  OAI2BB1X1 U23 ( .A0N(\u_div/PartRem[9][2] ), .A1N(n46), .B0(n11), .Y(n67) );
  MXI2X1 U24 ( .A(\u_div/PartRem[10][2] ), .B(\u_div/SumTmp[9][2] ), .S0(n66), 
        .Y(n11) );
  OAI2BB1X1 U25 ( .A0N(\u_div/PartRem[8][2] ), .A1N(n45), .B0(n12), .Y(n68) );
  MXI2X1 U26 ( .A(\u_div/PartRem[9][2] ), .B(\u_div/SumTmp[8][2] ), .S0(n67), 
        .Y(n12) );
  OAI2BB1X1 U27 ( .A0N(\u_div/PartRem[7][2] ), .A1N(n44), .B0(n13), .Y(n69) );
  MXI2X1 U28 ( .A(\u_div/PartRem[8][2] ), .B(\u_div/SumTmp[7][2] ), .S0(n68), 
        .Y(n13) );
  OAI2BB1X1 U29 ( .A0N(\u_div/PartRem[6][2] ), .A1N(n43), .B0(n14), .Y(n70) );
  MXI2X1 U30 ( .A(\u_div/PartRem[7][2] ), .B(\u_div/SumTmp[6][2] ), .S0(n69), 
        .Y(n14) );
  OAI2BB1X1 U31 ( .A0N(\u_div/PartRem[5][2] ), .A1N(n42), .B0(n15), .Y(n71) );
  MXI2X1 U32 ( .A(\u_div/PartRem[6][2] ), .B(\u_div/SumTmp[5][2] ), .S0(n70), 
        .Y(n15) );
  OAI2BB1X1 U33 ( .A0N(\u_div/PartRem[4][2] ), .A1N(n41), .B0(n16), .Y(n72) );
  MXI2X1 U34 ( .A(\u_div/PartRem[5][2] ), .B(\u_div/SumTmp[4][2] ), .S0(n71), 
        .Y(n16) );
  OAI2BB1X1 U35 ( .A0N(\u_div/PartRem[3][2] ), .A1N(n40), .B0(n17), .Y(n73) );
  MXI2X1 U36 ( .A(\u_div/PartRem[4][2] ), .B(\u_div/SumTmp[3][2] ), .S0(n72), 
        .Y(n17) );
  CLKINVX1 U37 ( .A(\u_div/CryTmp[3][1] ), .Y(n35) );
  CLKINVX1 U38 ( .A(\u_div/CryTmp[2][1] ), .Y(n36) );
  CLKINVX1 U39 ( .A(\u_div/CryTmp[1][1] ), .Y(n37) );
  INVXL U40 ( .A(\u_div/CryTmp[0][1] ), .Y(n19) );
  OAI2BB1X1 U41 ( .A0N(\u_div/PartRem[18][2] ), .A1N(n55), .B0(n18), .Y(n58)
         );
  MXI2X1 U42 ( .A(a[20]), .B(\u_div/SumTmp[18][2] ), .S0(n57), .Y(n18) );
  CLKINVX1 U43 ( .A(\u_div/CryTmp[18][1] ), .Y(n20) );
  CLKINVX1 U44 ( .A(\u_div/CryTmp[17][1] ), .Y(n21) );
  CLKINVX1 U45 ( .A(\u_div/CryTmp[16][1] ), .Y(n22) );
  CLKINVX1 U46 ( .A(\u_div/CryTmp[15][1] ), .Y(n23) );
  CLKINVX1 U47 ( .A(\u_div/CryTmp[14][1] ), .Y(n24) );
  CLKINVX1 U48 ( .A(\u_div/CryTmp[13][1] ), .Y(n25) );
  CLKINVX1 U49 ( .A(\u_div/CryTmp[12][1] ), .Y(n26) );
  CLKINVX1 U50 ( .A(\u_div/CryTmp[11][1] ), .Y(n27) );
  CLKINVX1 U51 ( .A(\u_div/CryTmp[10][1] ), .Y(n28) );
  CLKINVX1 U52 ( .A(\u_div/CryTmp[9][1] ), .Y(n29) );
  CLKINVX1 U53 ( .A(\u_div/CryTmp[8][1] ), .Y(n30) );
  CLKINVX1 U54 ( .A(\u_div/CryTmp[7][1] ), .Y(n31) );
  CLKINVX1 U55 ( .A(\u_div/CryTmp[6][1] ), .Y(n32) );
  CLKINVX1 U56 ( .A(\u_div/CryTmp[5][1] ), .Y(n33) );
  CLKINVX1 U57 ( .A(\u_div/CryTmp[4][1] ), .Y(n34) );
  XOR2X1 U58 ( .A(\u_div/PartRem[1][2] ), .B(n38), .Y(\u_div/SumTmp[0][2] ) );
  OR2X1 U59 ( .A(\u_div/CryTmp[1][1] ), .B(\u_div/PartRem[2][1] ), .Y(n39) );
  XNOR2X1 U60 ( .A(\u_div/PartRem[2][1] ), .B(\u_div/CryTmp[1][1] ), .Y(
        \u_div/SumTmp[1][1] ) );
  XOR2X1 U61 ( .A(\u_div/PartRem[2][2] ), .B(n39), .Y(\u_div/SumTmp[1][2] ) );
  OR2X1 U62 ( .A(\u_div/CryTmp[2][1] ), .B(\u_div/PartRem[3][1] ), .Y(n40) );
  XNOR2X1 U63 ( .A(\u_div/PartRem[3][1] ), .B(\u_div/CryTmp[2][1] ), .Y(
        \u_div/SumTmp[2][1] ) );
  XOR2X1 U64 ( .A(\u_div/PartRem[3][2] ), .B(n40), .Y(\u_div/SumTmp[2][2] ) );
  OR2X1 U65 ( .A(\u_div/CryTmp[3][1] ), .B(\u_div/PartRem[4][1] ), .Y(n41) );
  XNOR2X1 U66 ( .A(\u_div/PartRem[4][1] ), .B(\u_div/CryTmp[3][1] ), .Y(
        \u_div/SumTmp[3][1] ) );
  XOR2X1 U67 ( .A(\u_div/PartRem[4][2] ), .B(n41), .Y(\u_div/SumTmp[3][2] ) );
  OR2X1 U68 ( .A(\u_div/CryTmp[4][1] ), .B(\u_div/PartRem[5][1] ), .Y(n42) );
  XNOR2X1 U69 ( .A(\u_div/PartRem[5][1] ), .B(\u_div/CryTmp[4][1] ), .Y(
        \u_div/SumTmp[4][1] ) );
  XOR2X1 U70 ( .A(\u_div/PartRem[5][2] ), .B(n42), .Y(\u_div/SumTmp[4][2] ) );
  OR2X1 U71 ( .A(\u_div/CryTmp[5][1] ), .B(\u_div/PartRem[6][1] ), .Y(n43) );
  XNOR2X1 U72 ( .A(\u_div/PartRem[6][1] ), .B(\u_div/CryTmp[5][1] ), .Y(
        \u_div/SumTmp[5][1] ) );
  XOR2X1 U73 ( .A(\u_div/PartRem[6][2] ), .B(n43), .Y(\u_div/SumTmp[5][2] ) );
  OR2X1 U74 ( .A(\u_div/CryTmp[6][1] ), .B(\u_div/PartRem[7][1] ), .Y(n44) );
  XNOR2X1 U75 ( .A(\u_div/PartRem[7][1] ), .B(\u_div/CryTmp[6][1] ), .Y(
        \u_div/SumTmp[6][1] ) );
  XOR2X1 U76 ( .A(\u_div/PartRem[7][2] ), .B(n44), .Y(\u_div/SumTmp[6][2] ) );
  OR2X1 U77 ( .A(\u_div/CryTmp[7][1] ), .B(\u_div/PartRem[8][1] ), .Y(n45) );
  XNOR2X1 U78 ( .A(\u_div/PartRem[8][1] ), .B(\u_div/CryTmp[7][1] ), .Y(
        \u_div/SumTmp[7][1] ) );
  XOR2X1 U79 ( .A(\u_div/PartRem[8][2] ), .B(n45), .Y(\u_div/SumTmp[7][2] ) );
  OR2X1 U80 ( .A(\u_div/CryTmp[8][1] ), .B(\u_div/PartRem[9][1] ), .Y(n46) );
  XNOR2X1 U81 ( .A(\u_div/PartRem[9][1] ), .B(\u_div/CryTmp[8][1] ), .Y(
        \u_div/SumTmp[8][1] ) );
  XOR2X1 U82 ( .A(\u_div/PartRem[9][2] ), .B(n46), .Y(\u_div/SumTmp[8][2] ) );
  OR2X1 U83 ( .A(\u_div/CryTmp[9][1] ), .B(\u_div/PartRem[10][1] ), .Y(n47) );
  XNOR2X1 U84 ( .A(\u_div/PartRem[10][1] ), .B(\u_div/CryTmp[9][1] ), .Y(
        \u_div/SumTmp[9][1] ) );
  XOR2X1 U85 ( .A(\u_div/PartRem[10][2] ), .B(n47), .Y(\u_div/SumTmp[9][2] )
         );
  OR2X1 U86 ( .A(\u_div/CryTmp[10][1] ), .B(\u_div/PartRem[11][1] ), .Y(n48)
         );
  XNOR2X1 U87 ( .A(\u_div/PartRem[11][1] ), .B(\u_div/CryTmp[10][1] ), .Y(
        \u_div/SumTmp[10][1] ) );
  XOR2X1 U88 ( .A(\u_div/PartRem[11][2] ), .B(n48), .Y(\u_div/SumTmp[10][2] )
         );
  OR2X1 U89 ( .A(\u_div/CryTmp[11][1] ), .B(\u_div/PartRem[12][1] ), .Y(n49)
         );
  XNOR2X1 U90 ( .A(\u_div/PartRem[12][1] ), .B(\u_div/CryTmp[11][1] ), .Y(
        \u_div/SumTmp[11][1] ) );
  XOR2X1 U91 ( .A(\u_div/PartRem[12][2] ), .B(n49), .Y(\u_div/SumTmp[11][2] )
         );
  OR2X1 U92 ( .A(\u_div/CryTmp[12][1] ), .B(\u_div/PartRem[13][1] ), .Y(n50)
         );
  XNOR2X1 U93 ( .A(\u_div/PartRem[13][1] ), .B(\u_div/CryTmp[12][1] ), .Y(
        \u_div/SumTmp[12][1] ) );
  XOR2X1 U94 ( .A(\u_div/PartRem[13][2] ), .B(n50), .Y(\u_div/SumTmp[12][2] )
         );
  OR2X1 U95 ( .A(\u_div/CryTmp[13][1] ), .B(\u_div/PartRem[14][1] ), .Y(n51)
         );
  XNOR2X1 U96 ( .A(\u_div/PartRem[14][1] ), .B(\u_div/CryTmp[13][1] ), .Y(
        \u_div/SumTmp[13][1] ) );
  XOR2X1 U97 ( .A(\u_div/PartRem[14][2] ), .B(n51), .Y(\u_div/SumTmp[13][2] )
         );
  OR2X1 U98 ( .A(\u_div/CryTmp[14][1] ), .B(\u_div/PartRem[15][1] ), .Y(n52)
         );
  XNOR2X1 U99 ( .A(\u_div/PartRem[15][1] ), .B(\u_div/CryTmp[14][1] ), .Y(
        \u_div/SumTmp[14][1] ) );
  XOR2X1 U100 ( .A(\u_div/PartRem[15][2] ), .B(n52), .Y(\u_div/SumTmp[14][2] )
         );
  OR2X1 U101 ( .A(\u_div/CryTmp[15][1] ), .B(\u_div/PartRem[16][1] ), .Y(n53)
         );
  XNOR2X1 U102 ( .A(\u_div/PartRem[16][1] ), .B(\u_div/CryTmp[15][1] ), .Y(
        \u_div/SumTmp[15][1] ) );
  XOR2X1 U103 ( .A(\u_div/PartRem[16][2] ), .B(n53), .Y(\u_div/SumTmp[15][2] )
         );
  OR2X1 U104 ( .A(\u_div/CryTmp[16][1] ), .B(\u_div/PartRem[17][1] ), .Y(n54)
         );
  XNOR2X1 U105 ( .A(\u_div/PartRem[17][1] ), .B(\u_div/CryTmp[16][1] ), .Y(
        \u_div/SumTmp[16][1] ) );
  XOR2X1 U106 ( .A(\u_div/PartRem[17][2] ), .B(n54), .Y(\u_div/SumTmp[16][2] )
         );
  OR2X1 U107 ( .A(\u_div/CryTmp[17][1] ), .B(\u_div/PartRem[18][1] ), .Y(n55)
         );
  XNOR2X1 U108 ( .A(\u_div/PartRem[18][1] ), .B(\u_div/CryTmp[17][1] ), .Y(
        \u_div/SumTmp[17][1] ) );
  XOR2X1 U109 ( .A(\u_div/PartRem[18][2] ), .B(n55), .Y(\u_div/SumTmp[17][2] )
         );
  NOR2X1 U110 ( .A(\u_div/CryTmp[18][1] ), .B(\u_div/CryTmp[19][1] ), .Y(n56)
         );
  NOR2BX1 U111 ( .AN(a[20]), .B(n56), .Y(n57) );
  XNOR2X1 U112 ( .A(\u_div/CryTmp[19][1] ), .B(\u_div/CryTmp[18][1] ), .Y(
        \u_div/SumTmp[18][1] ) );
  XNOR2X1 U113 ( .A(a[20]), .B(n56), .Y(\u_div/SumTmp[18][2] ) );
endmodule


module CONT_DW_div_uns_15 ( a, b, quotient, remainder, divide_by_0 );
  input [20:0] a;
  input [2:0] b;
  output [20:0] quotient;
  output [2:0] remainder;
  output divide_by_0;
  wire   n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, \u_div/SumTmp[0][1] , \u_div/SumTmp[0][2] ,
         \u_div/SumTmp[1][1] , \u_div/SumTmp[1][2] , \u_div/SumTmp[2][1] ,
         \u_div/SumTmp[2][2] , \u_div/SumTmp[3][1] , \u_div/SumTmp[3][2] ,
         \u_div/SumTmp[4][1] , \u_div/SumTmp[4][2] , \u_div/SumTmp[5][1] ,
         \u_div/SumTmp[5][2] , \u_div/SumTmp[6][1] , \u_div/SumTmp[6][2] ,
         \u_div/SumTmp[7][1] , \u_div/SumTmp[7][2] , \u_div/SumTmp[8][1] ,
         \u_div/SumTmp[8][2] , \u_div/SumTmp[9][1] , \u_div/SumTmp[9][2] ,
         \u_div/SumTmp[10][1] , \u_div/SumTmp[10][2] , \u_div/SumTmp[11][1] ,
         \u_div/SumTmp[11][2] , \u_div/SumTmp[12][1] , \u_div/SumTmp[12][2] ,
         \u_div/SumTmp[13][1] , \u_div/SumTmp[13][2] , \u_div/SumTmp[14][1] ,
         \u_div/SumTmp[14][2] , \u_div/SumTmp[15][1] , \u_div/SumTmp[15][2] ,
         \u_div/SumTmp[16][1] , \u_div/SumTmp[16][2] , \u_div/SumTmp[17][1] ,
         \u_div/SumTmp[17][2] , \u_div/SumTmp[18][1] , \u_div/SumTmp[18][2] ,
         \u_div/CryTmp[0][1] , \u_div/CryTmp[1][1] , \u_div/CryTmp[2][1] ,
         \u_div/CryTmp[3][1] , \u_div/CryTmp[4][1] , \u_div/CryTmp[5][1] ,
         \u_div/CryTmp[6][1] , \u_div/CryTmp[7][1] , \u_div/CryTmp[8][1] ,
         \u_div/CryTmp[9][1] , \u_div/CryTmp[10][1] , \u_div/CryTmp[11][1] ,
         \u_div/CryTmp[12][1] , \u_div/CryTmp[13][1] , \u_div/CryTmp[14][1] ,
         \u_div/CryTmp[15][1] , \u_div/CryTmp[16][1] , \u_div/CryTmp[17][1] ,
         \u_div/CryTmp[18][1] , \u_div/CryTmp[19][1] , \u_div/PartRem[1][1] ,
         \u_div/PartRem[1][2] , \u_div/PartRem[2][1] , \u_div/PartRem[2][2] ,
         \u_div/PartRem[3][1] , \u_div/PartRem[3][2] , \u_div/PartRem[4][1] ,
         \u_div/PartRem[4][2] , \u_div/PartRem[5][1] , \u_div/PartRem[5][2] ,
         \u_div/PartRem[6][1] , \u_div/PartRem[6][2] , \u_div/PartRem[7][1] ,
         \u_div/PartRem[7][2] , \u_div/PartRem[8][1] , \u_div/PartRem[8][2] ,
         \u_div/PartRem[9][1] , \u_div/PartRem[9][2] , \u_div/PartRem[10][1] ,
         \u_div/PartRem[10][2] , \u_div/PartRem[11][1] ,
         \u_div/PartRem[11][2] , \u_div/PartRem[12][1] ,
         \u_div/PartRem[12][2] , \u_div/PartRem[13][1] ,
         \u_div/PartRem[13][2] , \u_div/PartRem[14][1] ,
         \u_div/PartRem[14][2] , \u_div/PartRem[15][1] ,
         \u_div/PartRem[15][2] , \u_div/PartRem[16][1] ,
         \u_div/PartRem[16][2] , \u_div/PartRem[17][1] ,
         \u_div/PartRem[17][2] , \u_div/PartRem[18][1] ,
         \u_div/PartRem[18][2] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56;
  assign \u_div/CryTmp[0][1]  = a[0];
  assign \u_div/CryTmp[1][1]  = a[1];
  assign \u_div/CryTmp[2][1]  = a[2];
  assign \u_div/CryTmp[3][1]  = a[3];
  assign \u_div/CryTmp[4][1]  = a[4];
  assign \u_div/CryTmp[5][1]  = a[5];
  assign \u_div/CryTmp[6][1]  = a[6];
  assign \u_div/CryTmp[7][1]  = a[7];
  assign \u_div/CryTmp[8][1]  = a[8];
  assign \u_div/CryTmp[9][1]  = a[9];
  assign \u_div/CryTmp[10][1]  = a[10];
  assign \u_div/CryTmp[11][1]  = a[11];
  assign \u_div/CryTmp[12][1]  = a[12];
  assign \u_div/CryTmp[13][1]  = a[13];
  assign \u_div/CryTmp[14][1]  = a[14];
  assign \u_div/CryTmp[15][1]  = a[15];
  assign \u_div/CryTmp[16][1]  = a[16];
  assign \u_div/CryTmp[17][1]  = a[17];
  assign \u_div/CryTmp[18][1]  = a[18];
  assign \u_div/CryTmp[19][1]  = a[19];

  CLKMX2X2 \u_div/u_mx_PartRem_0_4_1  ( .A(\u_div/PartRem[5][1] ), .B(
        \u_div/SumTmp[4][1] ), .S0(n71), .Y(\u_div/PartRem[4][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_5_1  ( .A(\u_div/PartRem[6][1] ), .B(
        \u_div/SumTmp[5][1] ), .S0(n70), .Y(\u_div/PartRem[5][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_6_1  ( .A(\u_div/PartRem[7][1] ), .B(
        \u_div/SumTmp[6][1] ), .S0(n69), .Y(\u_div/PartRem[6][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_7_1  ( .A(\u_div/PartRem[8][1] ), .B(
        \u_div/SumTmp[7][1] ), .S0(n68), .Y(\u_div/PartRem[7][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_8_1  ( .A(\u_div/PartRem[9][1] ), .B(
        \u_div/SumTmp[8][1] ), .S0(n67), .Y(\u_div/PartRem[8][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_9_1  ( .A(\u_div/PartRem[10][1] ), .B(
        \u_div/SumTmp[9][1] ), .S0(n66), .Y(\u_div/PartRem[9][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_10_1  ( .A(\u_div/PartRem[11][1] ), .B(
        \u_div/SumTmp[10][1] ), .S0(n65), .Y(\u_div/PartRem[10][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_11_1  ( .A(\u_div/PartRem[12][1] ), .B(
        \u_div/SumTmp[11][1] ), .S0(n64), .Y(\u_div/PartRem[11][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_12_1  ( .A(\u_div/PartRem[13][1] ), .B(
        \u_div/SumTmp[12][1] ), .S0(n63), .Y(\u_div/PartRem[12][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_13_1  ( .A(\u_div/PartRem[14][1] ), .B(
        \u_div/SumTmp[13][1] ), .S0(n62), .Y(\u_div/PartRem[13][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_14_1  ( .A(\u_div/PartRem[15][1] ), .B(
        \u_div/SumTmp[14][1] ), .S0(n61), .Y(\u_div/PartRem[14][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_15_1  ( .A(\u_div/PartRem[16][1] ), .B(
        \u_div/SumTmp[15][1] ), .S0(n60), .Y(\u_div/PartRem[15][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_16_1  ( .A(\u_div/PartRem[17][1] ), .B(
        \u_div/SumTmp[16][1] ), .S0(n59), .Y(\u_div/PartRem[16][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_17_1  ( .A(\u_div/PartRem[18][1] ), .B(
        \u_div/SumTmp[17][1] ), .S0(n58), .Y(\u_div/PartRem[17][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_18_1  ( .A(\u_div/CryTmp[19][1] ), .B(
        \u_div/SumTmp[18][1] ), .S0(n57), .Y(\u_div/PartRem[18][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_4_0  ( .A(\u_div/CryTmp[4][1] ), .B(n34), 
        .S0(n71), .Y(\u_div/PartRem[4][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_5_0  ( .A(\u_div/CryTmp[5][1] ), .B(n33), 
        .S0(n70), .Y(\u_div/PartRem[5][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_6_0  ( .A(\u_div/CryTmp[6][1] ), .B(n32), 
        .S0(n69), .Y(\u_div/PartRem[6][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_7_0  ( .A(\u_div/CryTmp[7][1] ), .B(n31), 
        .S0(n68), .Y(\u_div/PartRem[7][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_8_0  ( .A(\u_div/CryTmp[8][1] ), .B(n30), 
        .S0(n67), .Y(\u_div/PartRem[8][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_9_0  ( .A(\u_div/CryTmp[9][1] ), .B(n29), 
        .S0(n66), .Y(\u_div/PartRem[9][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_10_0  ( .A(\u_div/CryTmp[10][1] ), .B(n28), 
        .S0(n65), .Y(\u_div/PartRem[10][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_11_0  ( .A(\u_div/CryTmp[11][1] ), .B(n27), 
        .S0(n64), .Y(\u_div/PartRem[11][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_12_0  ( .A(\u_div/CryTmp[12][1] ), .B(n26), 
        .S0(n63), .Y(\u_div/PartRem[12][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_13_0  ( .A(\u_div/CryTmp[13][1] ), .B(n25), 
        .S0(n62), .Y(\u_div/PartRem[13][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_14_0  ( .A(\u_div/CryTmp[14][1] ), .B(n24), 
        .S0(n61), .Y(\u_div/PartRem[14][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_15_0  ( .A(\u_div/CryTmp[15][1] ), .B(n23), 
        .S0(n60), .Y(\u_div/PartRem[15][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_16_0  ( .A(\u_div/CryTmp[16][1] ), .B(n22), 
        .S0(n59), .Y(\u_div/PartRem[16][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_17_0  ( .A(\u_div/CryTmp[17][1] ), .B(n21), 
        .S0(n58), .Y(\u_div/PartRem[17][1] ) );
  MX2X1 \u_div/u_mx_PartRem_0_18_0  ( .A(\u_div/CryTmp[18][1] ), .B(n20), .S0(
        n57), .Y(\u_div/PartRem[18][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_1_1  ( .A(\u_div/PartRem[2][1] ), .B(
        \u_div/SumTmp[1][1] ), .S0(n74), .Y(\u_div/PartRem[1][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_2_1  ( .A(\u_div/PartRem[3][1] ), .B(
        \u_div/SumTmp[2][1] ), .S0(n73), .Y(\u_div/PartRem[2][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_3_1  ( .A(\u_div/PartRem[4][1] ), .B(
        \u_div/SumTmp[3][1] ), .S0(n72), .Y(\u_div/PartRem[3][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_1_0  ( .A(\u_div/CryTmp[1][1] ), .B(n37), 
        .S0(n74), .Y(\u_div/PartRem[1][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_2_0  ( .A(\u_div/CryTmp[2][1] ), .B(n36), 
        .S0(n73), .Y(\u_div/PartRem[2][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_3_0  ( .A(\u_div/CryTmp[3][1] ), .B(n35), 
        .S0(n72), .Y(\u_div/PartRem[3][1] ) );
  MX2XL \u_div/u_mx_PartRem_0_0_0  ( .A(\u_div/CryTmp[0][1] ), .B(n19), .S0(
        n75), .Y(remainder[0]) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_0_1  ( .A(\u_div/PartRem[1][1] ), .B(
        \u_div/SumTmp[0][1] ), .S0(n75), .Y(remainder[1]) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_0_2  ( .A(\u_div/PartRem[1][2] ), .B(
        \u_div/SumTmp[0][2] ), .S0(n75), .Y(remainder[2]) );
  OR2XL U1 ( .A(\u_div/CryTmp[0][1] ), .B(\u_div/PartRem[1][1] ), .Y(n38) );
  XNOR2XL U2 ( .A(\u_div/PartRem[1][1] ), .B(\u_div/CryTmp[0][1] ), .Y(
        \u_div/SumTmp[0][1] ) );
  OAI2BB1X1 U3 ( .A0N(\u_div/PartRem[2][2] ), .A1N(n39), .B0(n1), .Y(n74) );
  MXI2X1 U4 ( .A(\u_div/PartRem[3][2] ), .B(\u_div/SumTmp[2][2] ), .S0(n73), 
        .Y(n1) );
  OAI2BB1X1 U5 ( .A0N(\u_div/PartRem[1][2] ), .A1N(n38), .B0(n2), .Y(n75) );
  MXI2X1 U6 ( .A(\u_div/PartRem[2][2] ), .B(\u_div/SumTmp[1][2] ), .S0(n74), 
        .Y(n2) );
  OAI2BB1X1 U7 ( .A0N(\u_div/PartRem[17][2] ), .A1N(n54), .B0(n3), .Y(n59) );
  MXI2X1 U8 ( .A(\u_div/PartRem[18][2] ), .B(\u_div/SumTmp[17][2] ), .S0(n58), 
        .Y(n3) );
  OAI2BB1X1 U9 ( .A0N(\u_div/PartRem[16][2] ), .A1N(n53), .B0(n4), .Y(n60) );
  MXI2X1 U10 ( .A(\u_div/PartRem[17][2] ), .B(\u_div/SumTmp[16][2] ), .S0(n59), 
        .Y(n4) );
  OAI2BB1X1 U11 ( .A0N(\u_div/PartRem[15][2] ), .A1N(n52), .B0(n5), .Y(n61) );
  MXI2X1 U12 ( .A(\u_div/PartRem[16][2] ), .B(\u_div/SumTmp[15][2] ), .S0(n60), 
        .Y(n5) );
  OAI2BB1X1 U13 ( .A0N(\u_div/PartRem[14][2] ), .A1N(n51), .B0(n6), .Y(n62) );
  MXI2X1 U14 ( .A(\u_div/PartRem[15][2] ), .B(\u_div/SumTmp[14][2] ), .S0(n61), 
        .Y(n6) );
  OAI2BB1X1 U15 ( .A0N(\u_div/PartRem[13][2] ), .A1N(n50), .B0(n7), .Y(n63) );
  MXI2X1 U16 ( .A(\u_div/PartRem[14][2] ), .B(\u_div/SumTmp[13][2] ), .S0(n62), 
        .Y(n7) );
  OAI2BB1X1 U17 ( .A0N(\u_div/PartRem[12][2] ), .A1N(n49), .B0(n8), .Y(n64) );
  MXI2X1 U18 ( .A(\u_div/PartRem[13][2] ), .B(\u_div/SumTmp[12][2] ), .S0(n63), 
        .Y(n8) );
  OAI2BB1X1 U19 ( .A0N(\u_div/PartRem[11][2] ), .A1N(n48), .B0(n9), .Y(n65) );
  MXI2X1 U20 ( .A(\u_div/PartRem[12][2] ), .B(\u_div/SumTmp[11][2] ), .S0(n64), 
        .Y(n9) );
  OAI2BB1X1 U21 ( .A0N(\u_div/PartRem[10][2] ), .A1N(n47), .B0(n10), .Y(n66)
         );
  MXI2X1 U22 ( .A(\u_div/PartRem[11][2] ), .B(\u_div/SumTmp[10][2] ), .S0(n65), 
        .Y(n10) );
  OAI2BB1X1 U23 ( .A0N(\u_div/PartRem[9][2] ), .A1N(n46), .B0(n11), .Y(n67) );
  MXI2X1 U24 ( .A(\u_div/PartRem[10][2] ), .B(\u_div/SumTmp[9][2] ), .S0(n66), 
        .Y(n11) );
  OAI2BB1X1 U25 ( .A0N(\u_div/PartRem[8][2] ), .A1N(n45), .B0(n12), .Y(n68) );
  MXI2X1 U26 ( .A(\u_div/PartRem[9][2] ), .B(\u_div/SumTmp[8][2] ), .S0(n67), 
        .Y(n12) );
  OAI2BB1X1 U27 ( .A0N(\u_div/PartRem[7][2] ), .A1N(n44), .B0(n13), .Y(n69) );
  MXI2X1 U28 ( .A(\u_div/PartRem[8][2] ), .B(\u_div/SumTmp[7][2] ), .S0(n68), 
        .Y(n13) );
  OAI2BB1X1 U29 ( .A0N(\u_div/PartRem[6][2] ), .A1N(n43), .B0(n14), .Y(n70) );
  MXI2X1 U30 ( .A(\u_div/PartRem[7][2] ), .B(\u_div/SumTmp[6][2] ), .S0(n69), 
        .Y(n14) );
  OAI2BB1X1 U31 ( .A0N(\u_div/PartRem[5][2] ), .A1N(n42), .B0(n15), .Y(n71) );
  MXI2X1 U32 ( .A(\u_div/PartRem[6][2] ), .B(\u_div/SumTmp[5][2] ), .S0(n70), 
        .Y(n15) );
  OAI2BB1X1 U33 ( .A0N(\u_div/PartRem[4][2] ), .A1N(n41), .B0(n16), .Y(n72) );
  MXI2X1 U34 ( .A(\u_div/PartRem[5][2] ), .B(\u_div/SumTmp[4][2] ), .S0(n71), 
        .Y(n16) );
  OAI2BB1X1 U35 ( .A0N(\u_div/PartRem[3][2] ), .A1N(n40), .B0(n17), .Y(n73) );
  MXI2X1 U36 ( .A(\u_div/PartRem[4][2] ), .B(\u_div/SumTmp[3][2] ), .S0(n72), 
        .Y(n17) );
  CLKINVX1 U37 ( .A(\u_div/CryTmp[3][1] ), .Y(n35) );
  CLKINVX1 U38 ( .A(\u_div/CryTmp[2][1] ), .Y(n36) );
  CLKINVX1 U39 ( .A(\u_div/CryTmp[1][1] ), .Y(n37) );
  INVXL U40 ( .A(\u_div/CryTmp[0][1] ), .Y(n19) );
  OAI2BB1X1 U41 ( .A0N(\u_div/PartRem[18][2] ), .A1N(n55), .B0(n18), .Y(n58)
         );
  MXI2X1 U42 ( .A(a[20]), .B(\u_div/SumTmp[18][2] ), .S0(n57), .Y(n18) );
  CLKINVX1 U43 ( .A(\u_div/CryTmp[18][1] ), .Y(n20) );
  CLKINVX1 U44 ( .A(\u_div/CryTmp[17][1] ), .Y(n21) );
  CLKINVX1 U45 ( .A(\u_div/CryTmp[16][1] ), .Y(n22) );
  CLKINVX1 U46 ( .A(\u_div/CryTmp[15][1] ), .Y(n23) );
  CLKINVX1 U47 ( .A(\u_div/CryTmp[14][1] ), .Y(n24) );
  CLKINVX1 U48 ( .A(\u_div/CryTmp[13][1] ), .Y(n25) );
  CLKINVX1 U49 ( .A(\u_div/CryTmp[12][1] ), .Y(n26) );
  CLKINVX1 U50 ( .A(\u_div/CryTmp[11][1] ), .Y(n27) );
  CLKINVX1 U51 ( .A(\u_div/CryTmp[10][1] ), .Y(n28) );
  CLKINVX1 U52 ( .A(\u_div/CryTmp[9][1] ), .Y(n29) );
  CLKINVX1 U53 ( .A(\u_div/CryTmp[8][1] ), .Y(n30) );
  CLKINVX1 U54 ( .A(\u_div/CryTmp[7][1] ), .Y(n31) );
  CLKINVX1 U55 ( .A(\u_div/CryTmp[6][1] ), .Y(n32) );
  CLKINVX1 U56 ( .A(\u_div/CryTmp[5][1] ), .Y(n33) );
  CLKINVX1 U57 ( .A(\u_div/CryTmp[4][1] ), .Y(n34) );
  XOR2X1 U58 ( .A(\u_div/PartRem[1][2] ), .B(n38), .Y(\u_div/SumTmp[0][2] ) );
  OR2X1 U59 ( .A(\u_div/CryTmp[1][1] ), .B(\u_div/PartRem[2][1] ), .Y(n39) );
  XNOR2X1 U60 ( .A(\u_div/PartRem[2][1] ), .B(\u_div/CryTmp[1][1] ), .Y(
        \u_div/SumTmp[1][1] ) );
  XOR2X1 U61 ( .A(\u_div/PartRem[2][2] ), .B(n39), .Y(\u_div/SumTmp[1][2] ) );
  OR2X1 U62 ( .A(\u_div/CryTmp[2][1] ), .B(\u_div/PartRem[3][1] ), .Y(n40) );
  XNOR2X1 U63 ( .A(\u_div/PartRem[3][1] ), .B(\u_div/CryTmp[2][1] ), .Y(
        \u_div/SumTmp[2][1] ) );
  XOR2X1 U64 ( .A(\u_div/PartRem[3][2] ), .B(n40), .Y(\u_div/SumTmp[2][2] ) );
  OR2X1 U65 ( .A(\u_div/CryTmp[3][1] ), .B(\u_div/PartRem[4][1] ), .Y(n41) );
  XNOR2X1 U66 ( .A(\u_div/PartRem[4][1] ), .B(\u_div/CryTmp[3][1] ), .Y(
        \u_div/SumTmp[3][1] ) );
  XOR2X1 U67 ( .A(\u_div/PartRem[4][2] ), .B(n41), .Y(\u_div/SumTmp[3][2] ) );
  OR2X1 U68 ( .A(\u_div/CryTmp[4][1] ), .B(\u_div/PartRem[5][1] ), .Y(n42) );
  XNOR2X1 U69 ( .A(\u_div/PartRem[5][1] ), .B(\u_div/CryTmp[4][1] ), .Y(
        \u_div/SumTmp[4][1] ) );
  XOR2X1 U70 ( .A(\u_div/PartRem[5][2] ), .B(n42), .Y(\u_div/SumTmp[4][2] ) );
  OR2X1 U71 ( .A(\u_div/CryTmp[5][1] ), .B(\u_div/PartRem[6][1] ), .Y(n43) );
  XNOR2X1 U72 ( .A(\u_div/PartRem[6][1] ), .B(\u_div/CryTmp[5][1] ), .Y(
        \u_div/SumTmp[5][1] ) );
  XOR2X1 U73 ( .A(\u_div/PartRem[6][2] ), .B(n43), .Y(\u_div/SumTmp[5][2] ) );
  OR2X1 U74 ( .A(\u_div/CryTmp[6][1] ), .B(\u_div/PartRem[7][1] ), .Y(n44) );
  XNOR2X1 U75 ( .A(\u_div/PartRem[7][1] ), .B(\u_div/CryTmp[6][1] ), .Y(
        \u_div/SumTmp[6][1] ) );
  XOR2X1 U76 ( .A(\u_div/PartRem[7][2] ), .B(n44), .Y(\u_div/SumTmp[6][2] ) );
  OR2X1 U77 ( .A(\u_div/CryTmp[7][1] ), .B(\u_div/PartRem[8][1] ), .Y(n45) );
  XNOR2X1 U78 ( .A(\u_div/PartRem[8][1] ), .B(\u_div/CryTmp[7][1] ), .Y(
        \u_div/SumTmp[7][1] ) );
  XOR2X1 U79 ( .A(\u_div/PartRem[8][2] ), .B(n45), .Y(\u_div/SumTmp[7][2] ) );
  OR2X1 U80 ( .A(\u_div/CryTmp[8][1] ), .B(\u_div/PartRem[9][1] ), .Y(n46) );
  XNOR2X1 U81 ( .A(\u_div/PartRem[9][1] ), .B(\u_div/CryTmp[8][1] ), .Y(
        \u_div/SumTmp[8][1] ) );
  XOR2X1 U82 ( .A(\u_div/PartRem[9][2] ), .B(n46), .Y(\u_div/SumTmp[8][2] ) );
  OR2X1 U83 ( .A(\u_div/CryTmp[9][1] ), .B(\u_div/PartRem[10][1] ), .Y(n47) );
  XNOR2X1 U84 ( .A(\u_div/PartRem[10][1] ), .B(\u_div/CryTmp[9][1] ), .Y(
        \u_div/SumTmp[9][1] ) );
  XOR2X1 U85 ( .A(\u_div/PartRem[10][2] ), .B(n47), .Y(\u_div/SumTmp[9][2] )
         );
  OR2X1 U86 ( .A(\u_div/CryTmp[10][1] ), .B(\u_div/PartRem[11][1] ), .Y(n48)
         );
  XNOR2X1 U87 ( .A(\u_div/PartRem[11][1] ), .B(\u_div/CryTmp[10][1] ), .Y(
        \u_div/SumTmp[10][1] ) );
  XOR2X1 U88 ( .A(\u_div/PartRem[11][2] ), .B(n48), .Y(\u_div/SumTmp[10][2] )
         );
  OR2X1 U89 ( .A(\u_div/CryTmp[11][1] ), .B(\u_div/PartRem[12][1] ), .Y(n49)
         );
  XNOR2X1 U90 ( .A(\u_div/PartRem[12][1] ), .B(\u_div/CryTmp[11][1] ), .Y(
        \u_div/SumTmp[11][1] ) );
  XOR2X1 U91 ( .A(\u_div/PartRem[12][2] ), .B(n49), .Y(\u_div/SumTmp[11][2] )
         );
  OR2X1 U92 ( .A(\u_div/CryTmp[12][1] ), .B(\u_div/PartRem[13][1] ), .Y(n50)
         );
  XNOR2X1 U93 ( .A(\u_div/PartRem[13][1] ), .B(\u_div/CryTmp[12][1] ), .Y(
        \u_div/SumTmp[12][1] ) );
  XOR2X1 U94 ( .A(\u_div/PartRem[13][2] ), .B(n50), .Y(\u_div/SumTmp[12][2] )
         );
  OR2X1 U95 ( .A(\u_div/CryTmp[13][1] ), .B(\u_div/PartRem[14][1] ), .Y(n51)
         );
  XNOR2X1 U96 ( .A(\u_div/PartRem[14][1] ), .B(\u_div/CryTmp[13][1] ), .Y(
        \u_div/SumTmp[13][1] ) );
  XOR2X1 U97 ( .A(\u_div/PartRem[14][2] ), .B(n51), .Y(\u_div/SumTmp[13][2] )
         );
  OR2X1 U98 ( .A(\u_div/CryTmp[14][1] ), .B(\u_div/PartRem[15][1] ), .Y(n52)
         );
  XNOR2X1 U99 ( .A(\u_div/PartRem[15][1] ), .B(\u_div/CryTmp[14][1] ), .Y(
        \u_div/SumTmp[14][1] ) );
  XOR2X1 U100 ( .A(\u_div/PartRem[15][2] ), .B(n52), .Y(\u_div/SumTmp[14][2] )
         );
  OR2X1 U101 ( .A(\u_div/CryTmp[15][1] ), .B(\u_div/PartRem[16][1] ), .Y(n53)
         );
  XNOR2X1 U102 ( .A(\u_div/PartRem[16][1] ), .B(\u_div/CryTmp[15][1] ), .Y(
        \u_div/SumTmp[15][1] ) );
  XOR2X1 U103 ( .A(\u_div/PartRem[16][2] ), .B(n53), .Y(\u_div/SumTmp[15][2] )
         );
  OR2X1 U104 ( .A(\u_div/CryTmp[16][1] ), .B(\u_div/PartRem[17][1] ), .Y(n54)
         );
  XNOR2X1 U105 ( .A(\u_div/PartRem[17][1] ), .B(\u_div/CryTmp[16][1] ), .Y(
        \u_div/SumTmp[16][1] ) );
  XOR2X1 U106 ( .A(\u_div/PartRem[17][2] ), .B(n54), .Y(\u_div/SumTmp[16][2] )
         );
  OR2X1 U107 ( .A(\u_div/CryTmp[17][1] ), .B(\u_div/PartRem[18][1] ), .Y(n55)
         );
  XNOR2X1 U108 ( .A(\u_div/PartRem[18][1] ), .B(\u_div/CryTmp[17][1] ), .Y(
        \u_div/SumTmp[17][1] ) );
  XOR2X1 U109 ( .A(\u_div/PartRem[18][2] ), .B(n55), .Y(\u_div/SumTmp[17][2] )
         );
  NOR2X1 U110 ( .A(\u_div/CryTmp[18][1] ), .B(\u_div/CryTmp[19][1] ), .Y(n56)
         );
  NOR2BX1 U111 ( .AN(a[20]), .B(n56), .Y(n57) );
  XNOR2X1 U112 ( .A(\u_div/CryTmp[19][1] ), .B(\u_div/CryTmp[18][1] ), .Y(
        \u_div/SumTmp[18][1] ) );
  XNOR2X1 U113 ( .A(a[20]), .B(n56), .Y(\u_div/SumTmp[18][2] ) );
endmodule


module CONT_DW_div_uns_16 ( a, b, quotient, remainder, divide_by_0 );
  input [31:0] a;
  input [2:0] b;
  output [31:0] quotient;
  output [2:0] remainder;
  output divide_by_0;
  wire   n86, \u_div/SumTmp[0][0] , \u_div/SumTmp[1][0] , \u_div/SumTmp[2][0] ,
         \u_div/SumTmp[3][0] , \u_div/SumTmp[4][0] , \u_div/SumTmp[5][0] ,
         \u_div/SumTmp[6][0] , \u_div/SumTmp[7][0] , \u_div/SumTmp[8][0] ,
         \u_div/SumTmp[9][0] , \u_div/SumTmp[10][0] , \u_div/SumTmp[11][0] ,
         \u_div/SumTmp[12][0] , \u_div/SumTmp[13][0] , \u_div/SumTmp[14][0] ,
         \u_div/SumTmp[15][0] , \u_div/SumTmp[16][0] , \u_div/SumTmp[17][0] ,
         \u_div/SumTmp[18][0] , \u_div/SumTmp[19][0] , n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85;
  assign \u_div/SumTmp[0][0]  = a[0];
  assign \u_div/SumTmp[1][0]  = a[1];
  assign \u_div/SumTmp[2][0]  = a[2];
  assign \u_div/SumTmp[3][0]  = a[3];
  assign \u_div/SumTmp[4][0]  = a[4];
  assign \u_div/SumTmp[5][0]  = a[5];
  assign \u_div/SumTmp[6][0]  = a[6];
  assign \u_div/SumTmp[7][0]  = a[7];
  assign \u_div/SumTmp[8][0]  = a[8];
  assign \u_div/SumTmp[9][0]  = a[9];
  assign \u_div/SumTmp[10][0]  = a[10];
  assign \u_div/SumTmp[11][0]  = a[11];
  assign \u_div/SumTmp[12][0]  = a[12];
  assign \u_div/SumTmp[13][0]  = a[13];
  assign \u_div/SumTmp[14][0]  = a[14];
  assign \u_div/SumTmp[15][0]  = a[15];
  assign \u_div/SumTmp[16][0]  = a[16];
  assign \u_div/SumTmp[17][0]  = a[17];
  assign \u_div/SumTmp[18][0]  = a[18];
  assign \u_div/SumTmp[19][0]  = a[19];

  MX2XL \u_div/u_mx_PartRem_0_0_0  ( .A(\u_div/SumTmp[0][0] ), .B(
        \u_div/SumTmp[0][0] ), .S0(n86), .Y(remainder[0]) );
  OA21X2 U1 ( .A0(n62), .A1(n63), .B0(n61), .Y(n65) );
  MXI2X1 U2 ( .A(n60), .B(n59), .S0(n58), .Y(n61) );
  OA21X2 U3 ( .A0(n42), .A1(n43), .B0(n41), .Y(n45) );
  MXI2X1 U4 ( .A(n40), .B(n39), .S0(n38), .Y(n41) );
  OA21X2 U5 ( .A0(n27), .A1(n28), .B0(n26), .Y(n30) );
  MXI2X1 U6 ( .A(n25), .B(n24), .S0(n23), .Y(n26) );
  OA21X2 U7 ( .A0(n57), .A1(n58), .B0(n56), .Y(n60) );
  MXI2X1 U8 ( .A(n55), .B(n54), .S0(n53), .Y(n56) );
  OA21X2 U9 ( .A0(n77), .A1(n78), .B0(n76), .Y(n80) );
  MXI2X1 U10 ( .A(n75), .B(n74), .S0(n73), .Y(n76) );
  OA21X2 U11 ( .A0(n12), .A1(n13), .B0(n11), .Y(n15) );
  MXI2X1 U12 ( .A(n10), .B(n9), .S0(n8), .Y(n11) );
  OA21X2 U13 ( .A0(n7), .A1(n8), .B0(n6), .Y(n10) );
  OA21X2 U14 ( .A0(n52), .A1(n53), .B0(n51), .Y(n55) );
  MXI2X1 U15 ( .A(n50), .B(n49), .S0(n48), .Y(n51) );
  OA21X2 U16 ( .A0(n37), .A1(n38), .B0(n36), .Y(n40) );
  MXI2X1 U17 ( .A(n35), .B(n34), .S0(n33), .Y(n36) );
  OA21X2 U18 ( .A0(n22), .A1(n23), .B0(n21), .Y(n25) );
  MXI2X1 U19 ( .A(n20), .B(n19), .S0(n18), .Y(n21) );
  OA21X2 U20 ( .A0(n72), .A1(n73), .B0(n71), .Y(n75) );
  MXI2X1 U21 ( .A(n70), .B(n69), .S0(n68), .Y(n71) );
  OA21X2 U22 ( .A0(n47), .A1(n48), .B0(n46), .Y(n50) );
  OA21X2 U23 ( .A0(n32), .A1(n33), .B0(n31), .Y(n35) );
  OA21X2 U24 ( .A0(n17), .A1(n18), .B0(n16), .Y(n20) );
  OA21X2 U25 ( .A0(n67), .A1(n68), .B0(n66), .Y(n70) );
  OAI21X1 U26 ( .A0(n84), .A1(n83), .B0(n81), .Y(n86) );
  XNOR2XL U27 ( .A(n84), .B(n86), .Y(remainder[1]) );
  MXI2XL U28 ( .A(n80), .B(n79), .S0(n78), .Y(n81) );
  NOR2XL U29 ( .A(n80), .B(n77), .Y(n79) );
  NOR2XL U30 ( .A(n75), .B(n72), .Y(n74) );
  MXI2XL U31 ( .A(n83), .B(n82), .S0(n86), .Y(remainder[2]) );
  NOR2XL U32 ( .A(n70), .B(n67), .Y(n69) );
  MXI2XL U33 ( .A(n65), .B(n64), .S0(n63), .Y(n66) );
  NOR2XL U34 ( .A(n65), .B(n62), .Y(n64) );
  NOR2XL U35 ( .A(n60), .B(n57), .Y(n59) );
  NOR2XL U36 ( .A(n55), .B(n52), .Y(n54) );
  NOR2XL U37 ( .A(n10), .B(n7), .Y(n9) );
  MXI2XL U38 ( .A(n15), .B(n14), .S0(n13), .Y(n16) );
  NOR2XL U39 ( .A(n15), .B(n12), .Y(n14) );
  NOR2XL U40 ( .A(n20), .B(n17), .Y(n19) );
  NOR2XL U41 ( .A(n25), .B(n22), .Y(n24) );
  MXI2XL U42 ( .A(n30), .B(n29), .S0(n28), .Y(n31) );
  NOR2XL U43 ( .A(n30), .B(n27), .Y(n29) );
  NOR2XL U44 ( .A(n35), .B(n32), .Y(n34) );
  NOR2XL U45 ( .A(n40), .B(n37), .Y(n39) );
  MXI2XL U46 ( .A(n45), .B(n44), .S0(n43), .Y(n46) );
  NOR2XL U47 ( .A(n45), .B(n42), .Y(n44) );
  NOR2XL U48 ( .A(n50), .B(n47), .Y(n49) );
  CLKINVX1 U49 ( .A(\u_div/SumTmp[18][0] ), .Y(n85) );
  CLKINVX1 U50 ( .A(\u_div/SumTmp[1][0] ), .Y(n84) );
  CLKINVX1 U51 ( .A(\u_div/SumTmp[2][0] ), .Y(n77) );
  CLKINVX1 U52 ( .A(\u_div/SumTmp[3][0] ), .Y(n72) );
  CLKINVX1 U53 ( .A(\u_div/SumTmp[4][0] ), .Y(n67) );
  CLKINVX1 U54 ( .A(\u_div/SumTmp[5][0] ), .Y(n62) );
  CLKINVX1 U55 ( .A(\u_div/SumTmp[6][0] ), .Y(n57) );
  CLKINVX1 U56 ( .A(\u_div/SumTmp[7][0] ), .Y(n52) );
  CLKINVX1 U57 ( .A(\u_div/SumTmp[8][0] ), .Y(n47) );
  CLKINVX1 U58 ( .A(\u_div/SumTmp[9][0] ), .Y(n42) );
  CLKINVX1 U59 ( .A(\u_div/SumTmp[10][0] ), .Y(n37) );
  CLKINVX1 U60 ( .A(\u_div/SumTmp[11][0] ), .Y(n32) );
  CLKINVX1 U61 ( .A(\u_div/SumTmp[12][0] ), .Y(n27) );
  CLKINVX1 U62 ( .A(\u_div/SumTmp[13][0] ), .Y(n22) );
  CLKINVX1 U63 ( .A(\u_div/SumTmp[14][0] ), .Y(n17) );
  CLKINVX1 U64 ( .A(\u_div/SumTmp[15][0] ), .Y(n12) );
  CLKINVX1 U65 ( .A(\u_div/SumTmp[16][0] ), .Y(n7) );
  CLKINVX1 U66 ( .A(\u_div/SumTmp[17][0] ), .Y(n2) );
  NAND2X1 U67 ( .A(\u_div/SumTmp[18][0] ), .B(\u_div/SumTmp[19][0] ), .Y(n1)
         );
  MXI2X1 U68 ( .A(n85), .B(\u_div/SumTmp[18][0] ), .S0(n1), .Y(n3) );
  AOI2BB2X1 U69 ( .B0(n1), .B1(\u_div/SumTmp[19][0] ), .A0N(n3), .A1N(n2), .Y(
        n5) );
  XNOR2X1 U70 ( .A(n2), .B(n5), .Y(n8) );
  NOR2X1 U71 ( .A(n5), .B(n2), .Y(n4) );
  MXI2X1 U72 ( .A(n5), .B(n4), .S0(n3), .Y(n6) );
  XNOR2X1 U73 ( .A(n7), .B(n10), .Y(n13) );
  XNOR2X1 U74 ( .A(n12), .B(n15), .Y(n18) );
  XNOR2X1 U75 ( .A(n17), .B(n20), .Y(n23) );
  XNOR2X1 U76 ( .A(n22), .B(n25), .Y(n28) );
  XNOR2X1 U77 ( .A(n27), .B(n30), .Y(n33) );
  XNOR2X1 U78 ( .A(n32), .B(n35), .Y(n38) );
  XNOR2X1 U79 ( .A(n37), .B(n40), .Y(n43) );
  XNOR2X1 U80 ( .A(n42), .B(n45), .Y(n48) );
  XNOR2X1 U81 ( .A(n47), .B(n50), .Y(n53) );
  XNOR2X1 U82 ( .A(n52), .B(n55), .Y(n58) );
  XNOR2X1 U83 ( .A(n57), .B(n60), .Y(n63) );
  XNOR2X1 U84 ( .A(n62), .B(n65), .Y(n68) );
  XNOR2X1 U85 ( .A(n67), .B(n70), .Y(n73) );
  XNOR2X1 U86 ( .A(n72), .B(n75), .Y(n78) );
  XNOR2X1 U87 ( .A(n77), .B(n80), .Y(n83) );
  NAND2X1 U88 ( .A(\u_div/SumTmp[1][0] ), .B(n83), .Y(n82) );
endmodule


module CONT_DW01_inc_2 ( A, SUM );
  input [19:0] A;
  output [19:0] SUM;

  wire   [19:2] carry;

  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  ADDHXL U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHXL U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHXL U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHXL U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  ADDHXL U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  ADDHXL U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  ADDHXL U1_1_18 ( .A(A[18]), .B(carry[18]), .CO(carry[19]), .S(SUM[18]) );
  ADDHXL U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  XOR2X1 U1 ( .A(carry[19]), .B(A[19]), .Y(SUM[19]) );
  CLKINVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module CONT_DW01_inc_3 ( A, SUM );
  input [20:0] A;
  output [20:0] SUM;

  wire   [20:2] carry;

  CMPR22X2 U1_1_19 ( .A(A[19]), .B(carry[19]), .CO(SUM[20]), .S(SUM[19]) );
  CMPR22X2 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  CMPR22X2 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  CMPR22X2 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  CMPR22X2 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  CMPR22X2 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  CMPR22X2 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  CMPR22X2 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  CMPR22X2 U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  CMPR22X2 U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  CMPR22X2 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  CMPR22X2 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  CMPR22X2 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  CMPR22X2 U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  CMPR22X2 U1_1_18 ( .A(A[18]), .B(carry[18]), .CO(carry[19]), .S(SUM[18]) );
  CMPR22X2 U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  CMPR22X2 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  CMPR22X2 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  CMPR22X2 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INVX3 U1 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module CONT_DW_div_uns_17 ( a, b, quotient, remainder, divide_by_0 );
  input [19:0] a;
  input [2:0] b;
  output [19:0] quotient;
  output [2:0] remainder;
  output divide_by_0;
  wire   n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, \u_div/SumTmp[0][1] , \u_div/SumTmp[0][2] ,
         \u_div/SumTmp[1][1] , \u_div/SumTmp[1][2] , \u_div/SumTmp[2][1] ,
         \u_div/SumTmp[2][2] , \u_div/SumTmp[3][1] , \u_div/SumTmp[3][2] ,
         \u_div/SumTmp[4][1] , \u_div/SumTmp[4][2] , \u_div/SumTmp[5][1] ,
         \u_div/SumTmp[5][2] , \u_div/SumTmp[6][1] , \u_div/SumTmp[6][2] ,
         \u_div/SumTmp[7][1] , \u_div/SumTmp[7][2] , \u_div/SumTmp[8][1] ,
         \u_div/SumTmp[8][2] , \u_div/SumTmp[9][1] , \u_div/SumTmp[9][2] ,
         \u_div/SumTmp[10][1] , \u_div/SumTmp[10][2] , \u_div/SumTmp[11][1] ,
         \u_div/SumTmp[11][2] , \u_div/SumTmp[12][1] , \u_div/SumTmp[12][2] ,
         \u_div/SumTmp[13][1] , \u_div/SumTmp[13][2] , \u_div/SumTmp[14][1] ,
         \u_div/SumTmp[14][2] , \u_div/SumTmp[15][1] , \u_div/SumTmp[15][2] ,
         \u_div/SumTmp[16][1] , \u_div/SumTmp[16][2] , \u_div/SumTmp[17][1] ,
         \u_div/SumTmp[17][2] , \u_div/CryTmp[0][1] , \u_div/CryTmp[1][1] ,
         \u_div/CryTmp[2][1] , \u_div/CryTmp[3][1] , \u_div/CryTmp[4][1] ,
         \u_div/CryTmp[5][1] , \u_div/CryTmp[6][1] , \u_div/CryTmp[7][1] ,
         \u_div/CryTmp[8][1] , \u_div/CryTmp[9][1] , \u_div/CryTmp[10][1] ,
         \u_div/CryTmp[11][1] , \u_div/CryTmp[12][1] , \u_div/CryTmp[13][1] ,
         \u_div/CryTmp[14][1] , \u_div/CryTmp[15][1] , \u_div/CryTmp[16][1] ,
         \u_div/CryTmp[17][1] , \u_div/CryTmp[18][1] , \u_div/PartRem[1][1] ,
         \u_div/PartRem[1][2] , \u_div/PartRem[2][1] , \u_div/PartRem[2][2] ,
         \u_div/PartRem[3][1] , \u_div/PartRem[3][2] , \u_div/PartRem[4][1] ,
         \u_div/PartRem[4][2] , \u_div/PartRem[5][1] , \u_div/PartRem[5][2] ,
         \u_div/PartRem[6][1] , \u_div/PartRem[6][2] , \u_div/PartRem[7][1] ,
         \u_div/PartRem[7][2] , \u_div/PartRem[8][1] , \u_div/PartRem[8][2] ,
         \u_div/PartRem[9][1] , \u_div/PartRem[9][2] , \u_div/PartRem[10][1] ,
         \u_div/PartRem[10][2] , \u_div/PartRem[11][1] ,
         \u_div/PartRem[11][2] , \u_div/PartRem[12][1] ,
         \u_div/PartRem[12][2] , \u_div/PartRem[13][1] ,
         \u_div/PartRem[13][2] , \u_div/PartRem[14][1] ,
         \u_div/PartRem[14][2] , \u_div/PartRem[15][1] ,
         \u_div/PartRem[15][2] , \u_div/PartRem[16][1] ,
         \u_div/PartRem[16][2] , \u_div/PartRem[17][1] ,
         \u_div/PartRem[17][2] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53;
  assign \u_div/CryTmp[0][1]  = a[0];
  assign \u_div/CryTmp[1][1]  = a[1];
  assign \u_div/CryTmp[2][1]  = a[2];
  assign \u_div/CryTmp[3][1]  = a[3];
  assign \u_div/CryTmp[4][1]  = a[4];
  assign \u_div/CryTmp[5][1]  = a[5];
  assign \u_div/CryTmp[6][1]  = a[6];
  assign \u_div/CryTmp[7][1]  = a[7];
  assign \u_div/CryTmp[8][1]  = a[8];
  assign \u_div/CryTmp[9][1]  = a[9];
  assign \u_div/CryTmp[10][1]  = a[10];
  assign \u_div/CryTmp[11][1]  = a[11];
  assign \u_div/CryTmp[12][1]  = a[12];
  assign \u_div/CryTmp[13][1]  = a[13];
  assign \u_div/CryTmp[14][1]  = a[14];
  assign \u_div/CryTmp[15][1]  = a[15];
  assign \u_div/CryTmp[16][1]  = a[16];
  assign \u_div/CryTmp[17][1]  = a[17];
  assign \u_div/CryTmp[18][1]  = a[18];

  CLKMX2X2 \u_div/u_mx_PartRem_0_4_1  ( .A(\u_div/PartRem[5][1] ), .B(
        \u_div/SumTmp[4][1] ), .S0(n67), .Y(\u_div/PartRem[4][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_5_1  ( .A(\u_div/PartRem[6][1] ), .B(
        \u_div/SumTmp[5][1] ), .S0(n66), .Y(\u_div/PartRem[5][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_6_1  ( .A(\u_div/PartRem[7][1] ), .B(
        \u_div/SumTmp[6][1] ), .S0(n65), .Y(\u_div/PartRem[6][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_7_1  ( .A(\u_div/PartRem[8][1] ), .B(
        \u_div/SumTmp[7][1] ), .S0(n64), .Y(\u_div/PartRem[7][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_8_1  ( .A(\u_div/PartRem[9][1] ), .B(
        \u_div/SumTmp[8][1] ), .S0(n63), .Y(\u_div/PartRem[8][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_9_1  ( .A(\u_div/PartRem[10][1] ), .B(
        \u_div/SumTmp[9][1] ), .S0(n62), .Y(\u_div/PartRem[9][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_10_1  ( .A(\u_div/PartRem[11][1] ), .B(
        \u_div/SumTmp[10][1] ), .S0(n61), .Y(\u_div/PartRem[10][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_11_1  ( .A(\u_div/PartRem[12][1] ), .B(
        \u_div/SumTmp[11][1] ), .S0(n60), .Y(\u_div/PartRem[11][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_12_1  ( .A(\u_div/PartRem[13][1] ), .B(
        \u_div/SumTmp[12][1] ), .S0(n59), .Y(\u_div/PartRem[12][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_13_1  ( .A(\u_div/PartRem[14][1] ), .B(
        \u_div/SumTmp[13][1] ), .S0(n58), .Y(\u_div/PartRem[13][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_14_1  ( .A(\u_div/PartRem[15][1] ), .B(
        \u_div/SumTmp[14][1] ), .S0(n57), .Y(\u_div/PartRem[14][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_15_1  ( .A(\u_div/PartRem[16][1] ), .B(
        \u_div/SumTmp[15][1] ), .S0(n56), .Y(\u_div/PartRem[15][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_16_1  ( .A(\u_div/PartRem[17][1] ), .B(
        \u_div/SumTmp[16][1] ), .S0(n55), .Y(\u_div/PartRem[16][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_4_0  ( .A(\u_div/CryTmp[4][1] ), .B(n24), 
        .S0(n67), .Y(\u_div/PartRem[4][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_5_0  ( .A(\u_div/CryTmp[5][1] ), .B(n23), 
        .S0(n66), .Y(\u_div/PartRem[5][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_6_0  ( .A(\u_div/CryTmp[6][1] ), .B(n22), 
        .S0(n65), .Y(\u_div/PartRem[6][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_7_0  ( .A(\u_div/CryTmp[7][1] ), .B(n21), 
        .S0(n64), .Y(\u_div/PartRem[7][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_8_0  ( .A(\u_div/CryTmp[8][1] ), .B(n20), 
        .S0(n63), .Y(\u_div/PartRem[8][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_9_0  ( .A(\u_div/CryTmp[9][1] ), .B(n19), 
        .S0(n62), .Y(\u_div/PartRem[9][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_10_0  ( .A(\u_div/CryTmp[10][1] ), .B(n35), 
        .S0(n61), .Y(\u_div/PartRem[10][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_11_0  ( .A(\u_div/CryTmp[11][1] ), .B(n34), 
        .S0(n60), .Y(\u_div/PartRem[11][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_12_0  ( .A(\u_div/CryTmp[12][1] ), .B(n33), 
        .S0(n59), .Y(\u_div/PartRem[12][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_13_0  ( .A(\u_div/CryTmp[13][1] ), .B(n32), 
        .S0(n58), .Y(\u_div/PartRem[13][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_14_0  ( .A(\u_div/CryTmp[14][1] ), .B(n31), 
        .S0(n57), .Y(\u_div/PartRem[14][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_15_0  ( .A(\u_div/CryTmp[15][1] ), .B(n30), 
        .S0(n56), .Y(\u_div/PartRem[15][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_16_0  ( .A(\u_div/CryTmp[16][1] ), .B(n29), 
        .S0(n55), .Y(\u_div/PartRem[16][1] ) );
  MX2X1 \u_div/u_mx_PartRem_0_17_1  ( .A(\u_div/CryTmp[18][1] ), .B(
        \u_div/SumTmp[17][1] ), .S0(n54), .Y(\u_div/PartRem[17][2] ) );
  MX2X1 \u_div/u_mx_PartRem_0_17_0  ( .A(\u_div/CryTmp[17][1] ), .B(n28), .S0(
        n54), .Y(\u_div/PartRem[17][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_1_1  ( .A(\u_div/PartRem[2][1] ), .B(
        \u_div/SumTmp[1][1] ), .S0(n70), .Y(\u_div/PartRem[1][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_2_1  ( .A(\u_div/PartRem[3][1] ), .B(
        \u_div/SumTmp[2][1] ), .S0(n69), .Y(\u_div/PartRem[2][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_3_1  ( .A(\u_div/PartRem[4][1] ), .B(
        \u_div/SumTmp[3][1] ), .S0(n68), .Y(\u_div/PartRem[3][2] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_1_0  ( .A(\u_div/CryTmp[1][1] ), .B(n27), 
        .S0(n70), .Y(\u_div/PartRem[1][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_2_0  ( .A(\u_div/CryTmp[2][1] ), .B(n26), 
        .S0(n69), .Y(\u_div/PartRem[2][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_3_0  ( .A(\u_div/CryTmp[3][1] ), .B(n25), 
        .S0(n68), .Y(\u_div/PartRem[3][1] ) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_0_1  ( .A(\u_div/PartRem[1][1] ), .B(
        \u_div/SumTmp[0][1] ), .S0(n71), .Y(remainder[1]) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_0_0  ( .A(\u_div/CryTmp[0][1] ), .B(n18), 
        .S0(n71), .Y(remainder[0]) );
  CLKMX2X2 \u_div/u_mx_PartRem_0_0_2  ( .A(\u_div/PartRem[1][2] ), .B(
        \u_div/SumTmp[0][2] ), .S0(n71), .Y(remainder[2]) );
  NOR2X1 U1 ( .A(\u_div/CryTmp[17][1] ), .B(\u_div/CryTmp[18][1] ), .Y(n53) );
  XNOR2XL U2 ( .A(\u_div/CryTmp[18][1] ), .B(\u_div/CryTmp[17][1] ), .Y(
        \u_div/SumTmp[17][1] ) );
  OAI2BB1X1 U3 ( .A0N(\u_div/PartRem[2][2] ), .A1N(n37), .B0(n1), .Y(n70) );
  MXI2X1 U4 ( .A(\u_div/PartRem[3][2] ), .B(\u_div/SumTmp[2][2] ), .S0(n69), 
        .Y(n1) );
  OAI2BB1X1 U5 ( .A0N(\u_div/PartRem[1][2] ), .A1N(n36), .B0(n2), .Y(n71) );
  MXI2X1 U6 ( .A(\u_div/PartRem[2][2] ), .B(\u_div/SumTmp[1][2] ), .S0(n70), 
        .Y(n2) );
  OAI2BB1X1 U7 ( .A0N(\u_div/PartRem[16][2] ), .A1N(n51), .B0(n3), .Y(n56) );
  MXI2X1 U8 ( .A(\u_div/PartRem[17][2] ), .B(\u_div/SumTmp[16][2] ), .S0(n55), 
        .Y(n3) );
  OAI2BB1X1 U9 ( .A0N(\u_div/PartRem[15][2] ), .A1N(n50), .B0(n4), .Y(n57) );
  MXI2X1 U10 ( .A(\u_div/PartRem[16][2] ), .B(\u_div/SumTmp[15][2] ), .S0(n56), 
        .Y(n4) );
  OAI2BB1X1 U11 ( .A0N(\u_div/PartRem[14][2] ), .A1N(n49), .B0(n5), .Y(n58) );
  MXI2X1 U12 ( .A(\u_div/PartRem[15][2] ), .B(\u_div/SumTmp[14][2] ), .S0(n57), 
        .Y(n5) );
  OAI2BB1X1 U13 ( .A0N(\u_div/PartRem[13][2] ), .A1N(n48), .B0(n6), .Y(n59) );
  MXI2X1 U14 ( .A(\u_div/PartRem[14][2] ), .B(\u_div/SumTmp[13][2] ), .S0(n58), 
        .Y(n6) );
  OAI2BB1X1 U15 ( .A0N(\u_div/PartRem[12][2] ), .A1N(n47), .B0(n7), .Y(n60) );
  MXI2X1 U16 ( .A(\u_div/PartRem[13][2] ), .B(\u_div/SumTmp[12][2] ), .S0(n59), 
        .Y(n7) );
  OAI2BB1X1 U17 ( .A0N(\u_div/PartRem[11][2] ), .A1N(n46), .B0(n8), .Y(n61) );
  MXI2X1 U18 ( .A(\u_div/PartRem[12][2] ), .B(\u_div/SumTmp[11][2] ), .S0(n60), 
        .Y(n8) );
  OAI2BB1X1 U19 ( .A0N(\u_div/PartRem[10][2] ), .A1N(n45), .B0(n9), .Y(n62) );
  MXI2X1 U20 ( .A(\u_div/PartRem[11][2] ), .B(\u_div/SumTmp[10][2] ), .S0(n61), 
        .Y(n9) );
  OAI2BB1X1 U21 ( .A0N(\u_div/PartRem[9][2] ), .A1N(n44), .B0(n10), .Y(n63) );
  MXI2X1 U22 ( .A(\u_div/PartRem[10][2] ), .B(\u_div/SumTmp[9][2] ), .S0(n62), 
        .Y(n10) );
  OAI2BB1X1 U23 ( .A0N(\u_div/PartRem[8][2] ), .A1N(n43), .B0(n11), .Y(n64) );
  MXI2X1 U24 ( .A(\u_div/PartRem[9][2] ), .B(\u_div/SumTmp[8][2] ), .S0(n63), 
        .Y(n11) );
  OAI2BB1X1 U25 ( .A0N(\u_div/PartRem[7][2] ), .A1N(n42), .B0(n12), .Y(n65) );
  MXI2X1 U26 ( .A(\u_div/PartRem[8][2] ), .B(\u_div/SumTmp[7][2] ), .S0(n64), 
        .Y(n12) );
  OAI2BB1X1 U27 ( .A0N(\u_div/PartRem[6][2] ), .A1N(n41), .B0(n13), .Y(n66) );
  MXI2X1 U28 ( .A(\u_div/PartRem[7][2] ), .B(\u_div/SumTmp[6][2] ), .S0(n65), 
        .Y(n13) );
  OAI2BB1X1 U29 ( .A0N(\u_div/PartRem[5][2] ), .A1N(n40), .B0(n14), .Y(n67) );
  MXI2X1 U30 ( .A(\u_div/PartRem[6][2] ), .B(\u_div/SumTmp[5][2] ), .S0(n66), 
        .Y(n14) );
  OAI2BB1X1 U31 ( .A0N(\u_div/PartRem[4][2] ), .A1N(n39), .B0(n15), .Y(n68) );
  MXI2X1 U32 ( .A(\u_div/PartRem[5][2] ), .B(\u_div/SumTmp[4][2] ), .S0(n67), 
        .Y(n15) );
  OAI2BB1X1 U33 ( .A0N(\u_div/PartRem[3][2] ), .A1N(n38), .B0(n16), .Y(n69) );
  MXI2X1 U34 ( .A(\u_div/PartRem[4][2] ), .B(\u_div/SumTmp[3][2] ), .S0(n68), 
        .Y(n16) );
  CLKINVX1 U35 ( .A(\u_div/CryTmp[3][1] ), .Y(n25) );
  CLKINVX1 U36 ( .A(\u_div/CryTmp[2][1] ), .Y(n26) );
  CLKINVX1 U37 ( .A(\u_div/CryTmp[1][1] ), .Y(n27) );
  CLKINVX1 U38 ( .A(\u_div/CryTmp[0][1] ), .Y(n18) );
  OAI2BB1X1 U39 ( .A0N(\u_div/PartRem[17][2] ), .A1N(n52), .B0(n17), .Y(n55)
         );
  MXI2X1 U40 ( .A(a[19]), .B(\u_div/SumTmp[17][2] ), .S0(n54), .Y(n17) );
  CLKINVX1 U41 ( .A(\u_div/CryTmp[17][1] ), .Y(n28) );
  CLKINVX1 U42 ( .A(\u_div/CryTmp[16][1] ), .Y(n29) );
  CLKINVX1 U43 ( .A(\u_div/CryTmp[15][1] ), .Y(n30) );
  CLKINVX1 U44 ( .A(\u_div/CryTmp[14][1] ), .Y(n31) );
  CLKINVX1 U45 ( .A(\u_div/CryTmp[13][1] ), .Y(n32) );
  CLKINVX1 U46 ( .A(\u_div/CryTmp[12][1] ), .Y(n33) );
  CLKINVX1 U47 ( .A(\u_div/CryTmp[11][1] ), .Y(n34) );
  CLKINVX1 U48 ( .A(\u_div/CryTmp[10][1] ), .Y(n35) );
  CLKINVX1 U49 ( .A(\u_div/CryTmp[9][1] ), .Y(n19) );
  CLKINVX1 U50 ( .A(\u_div/CryTmp[8][1] ), .Y(n20) );
  CLKINVX1 U51 ( .A(\u_div/CryTmp[7][1] ), .Y(n21) );
  CLKINVX1 U52 ( .A(\u_div/CryTmp[6][1] ), .Y(n22) );
  CLKINVX1 U53 ( .A(\u_div/CryTmp[5][1] ), .Y(n23) );
  CLKINVX1 U54 ( .A(\u_div/CryTmp[4][1] ), .Y(n24) );
  OR2X1 U55 ( .A(\u_div/CryTmp[0][1] ), .B(\u_div/PartRem[1][1] ), .Y(n36) );
  XNOR2X1 U56 ( .A(\u_div/PartRem[1][1] ), .B(\u_div/CryTmp[0][1] ), .Y(
        \u_div/SumTmp[0][1] ) );
  XOR2X1 U57 ( .A(\u_div/PartRem[1][2] ), .B(n36), .Y(\u_div/SumTmp[0][2] ) );
  OR2X1 U58 ( .A(\u_div/CryTmp[1][1] ), .B(\u_div/PartRem[2][1] ), .Y(n37) );
  XNOR2X1 U59 ( .A(\u_div/PartRem[2][1] ), .B(\u_div/CryTmp[1][1] ), .Y(
        \u_div/SumTmp[1][1] ) );
  XOR2X1 U60 ( .A(\u_div/PartRem[2][2] ), .B(n37), .Y(\u_div/SumTmp[1][2] ) );
  OR2X1 U61 ( .A(\u_div/CryTmp[2][1] ), .B(\u_div/PartRem[3][1] ), .Y(n38) );
  XNOR2X1 U62 ( .A(\u_div/PartRem[3][1] ), .B(\u_div/CryTmp[2][1] ), .Y(
        \u_div/SumTmp[2][1] ) );
  XOR2X1 U63 ( .A(\u_div/PartRem[3][2] ), .B(n38), .Y(\u_div/SumTmp[2][2] ) );
  OR2X1 U64 ( .A(\u_div/CryTmp[3][1] ), .B(\u_div/PartRem[4][1] ), .Y(n39) );
  XNOR2X1 U65 ( .A(\u_div/PartRem[4][1] ), .B(\u_div/CryTmp[3][1] ), .Y(
        \u_div/SumTmp[3][1] ) );
  XOR2X1 U66 ( .A(\u_div/PartRem[4][2] ), .B(n39), .Y(\u_div/SumTmp[3][2] ) );
  OR2X1 U67 ( .A(\u_div/CryTmp[4][1] ), .B(\u_div/PartRem[5][1] ), .Y(n40) );
  XNOR2X1 U68 ( .A(\u_div/PartRem[5][1] ), .B(\u_div/CryTmp[4][1] ), .Y(
        \u_div/SumTmp[4][1] ) );
  XOR2X1 U69 ( .A(\u_div/PartRem[5][2] ), .B(n40), .Y(\u_div/SumTmp[4][2] ) );
  OR2X1 U70 ( .A(\u_div/CryTmp[5][1] ), .B(\u_div/PartRem[6][1] ), .Y(n41) );
  XNOR2X1 U71 ( .A(\u_div/PartRem[6][1] ), .B(\u_div/CryTmp[5][1] ), .Y(
        \u_div/SumTmp[5][1] ) );
  XOR2X1 U72 ( .A(\u_div/PartRem[6][2] ), .B(n41), .Y(\u_div/SumTmp[5][2] ) );
  OR2X1 U73 ( .A(\u_div/CryTmp[6][1] ), .B(\u_div/PartRem[7][1] ), .Y(n42) );
  XNOR2X1 U74 ( .A(\u_div/PartRem[7][1] ), .B(\u_div/CryTmp[6][1] ), .Y(
        \u_div/SumTmp[6][1] ) );
  XOR2X1 U75 ( .A(\u_div/PartRem[7][2] ), .B(n42), .Y(\u_div/SumTmp[6][2] ) );
  OR2X1 U76 ( .A(\u_div/CryTmp[7][1] ), .B(\u_div/PartRem[8][1] ), .Y(n43) );
  XNOR2X1 U77 ( .A(\u_div/PartRem[8][1] ), .B(\u_div/CryTmp[7][1] ), .Y(
        \u_div/SumTmp[7][1] ) );
  XOR2X1 U78 ( .A(\u_div/PartRem[8][2] ), .B(n43), .Y(\u_div/SumTmp[7][2] ) );
  OR2X1 U79 ( .A(\u_div/CryTmp[8][1] ), .B(\u_div/PartRem[9][1] ), .Y(n44) );
  XNOR2X1 U80 ( .A(\u_div/PartRem[9][1] ), .B(\u_div/CryTmp[8][1] ), .Y(
        \u_div/SumTmp[8][1] ) );
  XOR2X1 U81 ( .A(\u_div/PartRem[9][2] ), .B(n44), .Y(\u_div/SumTmp[8][2] ) );
  OR2X1 U82 ( .A(\u_div/CryTmp[9][1] ), .B(\u_div/PartRem[10][1] ), .Y(n45) );
  XNOR2X1 U83 ( .A(\u_div/PartRem[10][1] ), .B(\u_div/CryTmp[9][1] ), .Y(
        \u_div/SumTmp[9][1] ) );
  XOR2X1 U84 ( .A(\u_div/PartRem[10][2] ), .B(n45), .Y(\u_div/SumTmp[9][2] )
         );
  OR2X1 U85 ( .A(\u_div/CryTmp[10][1] ), .B(\u_div/PartRem[11][1] ), .Y(n46)
         );
  XNOR2X1 U86 ( .A(\u_div/PartRem[11][1] ), .B(\u_div/CryTmp[10][1] ), .Y(
        \u_div/SumTmp[10][1] ) );
  XOR2X1 U87 ( .A(\u_div/PartRem[11][2] ), .B(n46), .Y(\u_div/SumTmp[10][2] )
         );
  OR2X1 U88 ( .A(\u_div/CryTmp[11][1] ), .B(\u_div/PartRem[12][1] ), .Y(n47)
         );
  XNOR2X1 U89 ( .A(\u_div/PartRem[12][1] ), .B(\u_div/CryTmp[11][1] ), .Y(
        \u_div/SumTmp[11][1] ) );
  XOR2X1 U90 ( .A(\u_div/PartRem[12][2] ), .B(n47), .Y(\u_div/SumTmp[11][2] )
         );
  OR2X1 U91 ( .A(\u_div/CryTmp[12][1] ), .B(\u_div/PartRem[13][1] ), .Y(n48)
         );
  XNOR2X1 U92 ( .A(\u_div/PartRem[13][1] ), .B(\u_div/CryTmp[12][1] ), .Y(
        \u_div/SumTmp[12][1] ) );
  XOR2X1 U93 ( .A(\u_div/PartRem[13][2] ), .B(n48), .Y(\u_div/SumTmp[12][2] )
         );
  OR2X1 U94 ( .A(\u_div/CryTmp[13][1] ), .B(\u_div/PartRem[14][1] ), .Y(n49)
         );
  XNOR2X1 U95 ( .A(\u_div/PartRem[14][1] ), .B(\u_div/CryTmp[13][1] ), .Y(
        \u_div/SumTmp[13][1] ) );
  XOR2X1 U96 ( .A(\u_div/PartRem[14][2] ), .B(n49), .Y(\u_div/SumTmp[13][2] )
         );
  OR2X1 U97 ( .A(\u_div/CryTmp[14][1] ), .B(\u_div/PartRem[15][1] ), .Y(n50)
         );
  XNOR2X1 U98 ( .A(\u_div/PartRem[15][1] ), .B(\u_div/CryTmp[14][1] ), .Y(
        \u_div/SumTmp[14][1] ) );
  XOR2X1 U99 ( .A(\u_div/PartRem[15][2] ), .B(n50), .Y(\u_div/SumTmp[14][2] )
         );
  OR2X1 U100 ( .A(\u_div/CryTmp[15][1] ), .B(\u_div/PartRem[16][1] ), .Y(n51)
         );
  XNOR2X1 U101 ( .A(\u_div/PartRem[16][1] ), .B(\u_div/CryTmp[15][1] ), .Y(
        \u_div/SumTmp[15][1] ) );
  XOR2X1 U102 ( .A(\u_div/PartRem[16][2] ), .B(n51), .Y(\u_div/SumTmp[15][2] )
         );
  OR2X1 U103 ( .A(\u_div/CryTmp[16][1] ), .B(\u_div/PartRem[17][1] ), .Y(n52)
         );
  XNOR2X1 U104 ( .A(\u_div/PartRem[17][1] ), .B(\u_div/CryTmp[16][1] ), .Y(
        \u_div/SumTmp[16][1] ) );
  XOR2X1 U105 ( .A(\u_div/PartRem[17][2] ), .B(n52), .Y(\u_div/SumTmp[16][2] )
         );
  NOR2BX1 U106 ( .AN(a[19]), .B(n53), .Y(n54) );
  XNOR2X1 U107 ( .A(a[19]), .B(n53), .Y(\u_div/SumTmp[17][2] ) );
endmodule


module CONT_DW_div_uns_18 ( a, b, quotient, remainder, divide_by_0 );
  input [31:0] a;
  input [2:0] b;
  output [31:0] quotient;
  output [2:0] remainder;
  output divide_by_0;
  wire   n86, \u_div/SumTmp[0][0] , \u_div/SumTmp[1][0] , \u_div/SumTmp[2][0] ,
         \u_div/SumTmp[3][0] , \u_div/SumTmp[4][0] , \u_div/SumTmp[5][0] ,
         \u_div/SumTmp[6][0] , \u_div/SumTmp[7][0] , \u_div/SumTmp[8][0] ,
         \u_div/SumTmp[9][0] , \u_div/SumTmp[10][0] , \u_div/SumTmp[11][0] ,
         \u_div/SumTmp[12][0] , \u_div/SumTmp[13][0] , \u_div/SumTmp[14][0] ,
         \u_div/SumTmp[15][0] , \u_div/SumTmp[16][0] , \u_div/SumTmp[17][0] ,
         \u_div/SumTmp[18][0] , \u_div/SumTmp[19][0] , n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85;
  assign \u_div/SumTmp[0][0]  = a[0];
  assign \u_div/SumTmp[1][0]  = a[1];
  assign \u_div/SumTmp[2][0]  = a[2];
  assign \u_div/SumTmp[3][0]  = a[3];
  assign \u_div/SumTmp[4][0]  = a[4];
  assign \u_div/SumTmp[5][0]  = a[5];
  assign \u_div/SumTmp[6][0]  = a[6];
  assign \u_div/SumTmp[7][0]  = a[7];
  assign \u_div/SumTmp[8][0]  = a[8];
  assign \u_div/SumTmp[9][0]  = a[9];
  assign \u_div/SumTmp[10][0]  = a[10];
  assign \u_div/SumTmp[11][0]  = a[11];
  assign \u_div/SumTmp[12][0]  = a[12];
  assign \u_div/SumTmp[13][0]  = a[13];
  assign \u_div/SumTmp[14][0]  = a[14];
  assign \u_div/SumTmp[15][0]  = a[15];
  assign \u_div/SumTmp[16][0]  = a[16];
  assign \u_div/SumTmp[17][0]  = a[17];
  assign \u_div/SumTmp[18][0]  = a[18];
  assign \u_div/SumTmp[19][0]  = a[19];

  MX2XL \u_div/u_mx_PartRem_0_0_0  ( .A(\u_div/SumTmp[0][0] ), .B(
        \u_div/SumTmp[0][0] ), .S0(n86), .Y(remainder[0]) );
  OA21X2 U1 ( .A0(n47), .A1(n48), .B0(n46), .Y(n50) );
  MXI2X1 U2 ( .A(n45), .B(n44), .S0(n43), .Y(n46) );
  OA21X2 U3 ( .A0(n42), .A1(n43), .B0(n41), .Y(n45) );
  MXI2X1 U4 ( .A(n40), .B(n39), .S0(n38), .Y(n41) );
  OA21X2 U5 ( .A0(n67), .A1(n68), .B0(n66), .Y(n70) );
  MXI2X1 U6 ( .A(n65), .B(n64), .S0(n63), .Y(n66) );
  OA21X2 U7 ( .A0(n27), .A1(n28), .B0(n26), .Y(n30) );
  MXI2X1 U8 ( .A(n25), .B(n24), .S0(n23), .Y(n26) );
  OA21X2 U9 ( .A0(n52), .A1(n53), .B0(n51), .Y(n55) );
  OA21X2 U10 ( .A0(n12), .A1(n13), .B0(n11), .Y(n15) );
  MXI2X1 U11 ( .A(n10), .B(n9), .S0(n8), .Y(n11) );
  OA21X2 U12 ( .A0(n77), .A1(n78), .B0(n76), .Y(n80) );
  MXI2X1 U13 ( .A(n75), .B(n74), .S0(n73), .Y(n76) );
  OA21X2 U14 ( .A0(n7), .A1(n8), .B0(n6), .Y(n10) );
  OA21X2 U15 ( .A0(n37), .A1(n38), .B0(n36), .Y(n40) );
  MXI2X1 U16 ( .A(n35), .B(n34), .S0(n33), .Y(n36) );
  OA21X2 U17 ( .A0(n22), .A1(n23), .B0(n21), .Y(n25) );
  MXI2X1 U18 ( .A(n20), .B(n19), .S0(n18), .Y(n21) );
  OA21X2 U19 ( .A0(n62), .A1(n63), .B0(n61), .Y(n65) );
  MXI2X1 U20 ( .A(n60), .B(n59), .S0(n58), .Y(n61) );
  OAI21X1 U21 ( .A0(n84), .A1(n83), .B0(n81), .Y(n86) );
  OA21X2 U22 ( .A0(n32), .A1(n33), .B0(n31), .Y(n35) );
  OA21X2 U23 ( .A0(n17), .A1(n18), .B0(n16), .Y(n20) );
  OA21X2 U24 ( .A0(n57), .A1(n58), .B0(n56), .Y(n60) );
  OA21X2 U25 ( .A0(n72), .A1(n73), .B0(n71), .Y(n75) );
  MXI2XL U26 ( .A(n80), .B(n79), .S0(n78), .Y(n81) );
  NOR2XL U27 ( .A(n80), .B(n77), .Y(n79) );
  NOR2XL U28 ( .A(n75), .B(n72), .Y(n74) );
  XNOR2XL U29 ( .A(n84), .B(n86), .Y(remainder[1]) );
  MXI2XL U30 ( .A(n83), .B(n82), .S0(n86), .Y(remainder[2]) );
  MXI2XL U31 ( .A(n70), .B(n69), .S0(n68), .Y(n71) );
  NOR2XL U32 ( .A(n70), .B(n67), .Y(n69) );
  NOR2XL U33 ( .A(n65), .B(n62), .Y(n64) );
  NOR2XL U34 ( .A(n60), .B(n57), .Y(n59) );
  MXI2XL U35 ( .A(n55), .B(n54), .S0(n53), .Y(n56) );
  NOR2XL U36 ( .A(n55), .B(n52), .Y(n54) );
  NOR2XL U37 ( .A(n10), .B(n7), .Y(n9) );
  MXI2XL U38 ( .A(n15), .B(n14), .S0(n13), .Y(n16) );
  NOR2XL U39 ( .A(n15), .B(n12), .Y(n14) );
  NOR2XL U40 ( .A(n20), .B(n17), .Y(n19) );
  NOR2XL U41 ( .A(n25), .B(n22), .Y(n24) );
  MXI2XL U42 ( .A(n30), .B(n29), .S0(n28), .Y(n31) );
  NOR2XL U43 ( .A(n30), .B(n27), .Y(n29) );
  NOR2XL U44 ( .A(n35), .B(n32), .Y(n34) );
  NOR2XL U45 ( .A(n40), .B(n37), .Y(n39) );
  NOR2XL U46 ( .A(n45), .B(n42), .Y(n44) );
  MXI2XL U47 ( .A(n50), .B(n49), .S0(n48), .Y(n51) );
  NOR2XL U48 ( .A(n50), .B(n47), .Y(n49) );
  CLKINVX1 U49 ( .A(\u_div/SumTmp[18][0] ), .Y(n85) );
  CLKINVX1 U50 ( .A(\u_div/SumTmp[1][0] ), .Y(n84) );
  CLKINVX1 U51 ( .A(\u_div/SumTmp[2][0] ), .Y(n77) );
  CLKINVX1 U52 ( .A(\u_div/SumTmp[3][0] ), .Y(n72) );
  CLKINVX1 U53 ( .A(\u_div/SumTmp[4][0] ), .Y(n67) );
  CLKINVX1 U54 ( .A(\u_div/SumTmp[5][0] ), .Y(n62) );
  CLKINVX1 U55 ( .A(\u_div/SumTmp[6][0] ), .Y(n57) );
  CLKINVX1 U56 ( .A(\u_div/SumTmp[7][0] ), .Y(n52) );
  CLKINVX1 U57 ( .A(\u_div/SumTmp[8][0] ), .Y(n47) );
  CLKINVX1 U58 ( .A(\u_div/SumTmp[9][0] ), .Y(n42) );
  CLKINVX1 U59 ( .A(\u_div/SumTmp[10][0] ), .Y(n37) );
  CLKINVX1 U60 ( .A(\u_div/SumTmp[11][0] ), .Y(n32) );
  CLKINVX1 U61 ( .A(\u_div/SumTmp[12][0] ), .Y(n27) );
  CLKINVX1 U62 ( .A(\u_div/SumTmp[13][0] ), .Y(n22) );
  CLKINVX1 U63 ( .A(\u_div/SumTmp[14][0] ), .Y(n17) );
  CLKINVX1 U64 ( .A(\u_div/SumTmp[15][0] ), .Y(n12) );
  CLKINVX1 U65 ( .A(\u_div/SumTmp[16][0] ), .Y(n7) );
  CLKINVX1 U66 ( .A(\u_div/SumTmp[17][0] ), .Y(n2) );
  NAND2X1 U67 ( .A(\u_div/SumTmp[18][0] ), .B(\u_div/SumTmp[19][0] ), .Y(n1)
         );
  MXI2X1 U68 ( .A(n85), .B(\u_div/SumTmp[18][0] ), .S0(n1), .Y(n3) );
  AOI2BB2X1 U69 ( .B0(n1), .B1(\u_div/SumTmp[19][0] ), .A0N(n3), .A1N(n2), .Y(
        n5) );
  XNOR2X1 U70 ( .A(n2), .B(n5), .Y(n8) );
  NOR2X1 U71 ( .A(n5), .B(n2), .Y(n4) );
  MXI2X1 U72 ( .A(n5), .B(n4), .S0(n3), .Y(n6) );
  XNOR2X1 U73 ( .A(n7), .B(n10), .Y(n13) );
  XNOR2X1 U74 ( .A(n12), .B(n15), .Y(n18) );
  XNOR2X1 U75 ( .A(n17), .B(n20), .Y(n23) );
  XNOR2X1 U76 ( .A(n22), .B(n25), .Y(n28) );
  XNOR2X1 U77 ( .A(n27), .B(n30), .Y(n33) );
  XNOR2X1 U78 ( .A(n32), .B(n35), .Y(n38) );
  XNOR2X1 U79 ( .A(n37), .B(n40), .Y(n43) );
  XNOR2X1 U80 ( .A(n42), .B(n45), .Y(n48) );
  XNOR2X1 U81 ( .A(n47), .B(n50), .Y(n53) );
  XNOR2X1 U82 ( .A(n52), .B(n55), .Y(n58) );
  XNOR2X1 U83 ( .A(n57), .B(n60), .Y(n63) );
  XNOR2X1 U84 ( .A(n62), .B(n65), .Y(n68) );
  XNOR2X1 U85 ( .A(n67), .B(n70), .Y(n73) );
  XNOR2X1 U86 ( .A(n72), .B(n75), .Y(n78) );
  XNOR2X1 U87 ( .A(n77), .B(n80), .Y(n83) );
  NAND2X1 U88 ( .A(\u_div/SumTmp[1][0] ), .B(n83), .Y(n82) );
endmodule


module CONT_DW01_inc_4 ( A, SUM );
  input [19:0] A;
  output [19:0] SUM;

  wire   [19:2] carry;

  ADDHXL U1_1_18 ( .A(A[18]), .B(carry[18]), .CO(carry[19]), .S(SUM[18]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  ADDHXL U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  ADDHXL U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  ADDHXL U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  ADDHXL U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  ADDHXL U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADDHXL U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHXL U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHXL U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHXL U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(carry[19]), .B(A[19]), .Y(SUM[19]) );
  CLKINVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module CONT_DW_div_uns_19 ( a, b, quotient, remainder, divide_by_0 );
  input [31:0] a;
  input [3:0] b;
  output [31:0] quotient;
  output [3:0] remainder;
  output divide_by_0;
  wire   n130, \u_div/SumTmp[0][0] , \u_div/SumTmp[1][0] ,
         \u_div/SumTmp[2][0] , \u_div/SumTmp[3][0] , \u_div/SumTmp[4][0] ,
         \u_div/SumTmp[5][0] , \u_div/SumTmp[6][0] , \u_div/SumTmp[7][0] ,
         \u_div/SumTmp[8][0] , \u_div/SumTmp[9][0] , \u_div/SumTmp[10][0] ,
         \u_div/SumTmp[11][0] , \u_div/SumTmp[12][0] , \u_div/SumTmp[13][0] ,
         \u_div/SumTmp[14][0] , \u_div/SumTmp[15][0] , \u_div/SumTmp[16][0] ,
         \u_div/SumTmp[16][2] , \u_div/SumTmp[17][0] , \u_div/SumTmp[18][0] ,
         \u_div/SumTmp[19][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129;
  assign \u_div/SumTmp[0][0]  = a[0];
  assign \u_div/SumTmp[1][0]  = a[1];
  assign \u_div/SumTmp[2][0]  = a[2];
  assign \u_div/SumTmp[3][0]  = a[3];
  assign \u_div/SumTmp[4][0]  = a[4];
  assign \u_div/SumTmp[5][0]  = a[5];
  assign \u_div/SumTmp[6][0]  = a[6];
  assign \u_div/SumTmp[7][0]  = a[7];
  assign \u_div/SumTmp[8][0]  = a[8];
  assign \u_div/SumTmp[9][0]  = a[9];
  assign \u_div/SumTmp[10][0]  = a[10];
  assign \u_div/SumTmp[11][0]  = a[11];
  assign \u_div/SumTmp[12][0]  = a[12];
  assign \u_div/SumTmp[13][0]  = a[13];
  assign \u_div/SumTmp[14][0]  = a[14];
  assign \u_div/SumTmp[15][0]  = a[15];
  assign \u_div/SumTmp[16][0]  = a[16];
  assign \u_div/SumTmp[17][0]  = a[17];
  assign \u_div/SumTmp[18][0]  = a[18];
  assign \u_div/SumTmp[19][0]  = a[19];

  MX2XL \u_div/u_mx_PartRem_0_0_0  ( .A(\u_div/SumTmp[0][0] ), .B(
        \u_div/SumTmp[0][0] ), .S0(n130), .Y(remainder[0]) );
  OA21X2 U1 ( .A0(n100), .A1(n101), .B0(n97), .Y(n102) );
  AOI2BB2X2 U2 ( .B0(n1), .B1(\u_div/SumTmp[19][0] ), .A0N(n4), .A1N(n5), .Y(
        n6) );
  OA21X2 U3 ( .A0(n76), .A1(n77), .B0(n73), .Y(n78) );
  OA21X2 U4 ( .A0(n52), .A1(n53), .B0(n49), .Y(n54) );
  OA21X2 U5 ( .A0(n28), .A1(n29), .B0(n25), .Y(n30) );
  OA21X2 U6 ( .A0(n108), .A1(n109), .B0(n105), .Y(n110) );
  OA21X2 U7 ( .A0(n12), .A1(n13), .B0(n9), .Y(n14) );
  OA21X2 U8 ( .A0(n84), .A1(n85), .B0(n81), .Y(n86) );
  OA21X2 U9 ( .A0(n60), .A1(n61), .B0(n57), .Y(n62) );
  OA21X2 U10 ( .A0(n36), .A1(n37), .B0(n33), .Y(n38) );
  MXI2X2 U11 ( .A(n115), .B(n114), .S0(n118), .Y(n124) );
  OA21X2 U12 ( .A0(n92), .A1(n93), .B0(n89), .Y(n94) );
  OA21X2 U13 ( .A0(n68), .A1(n69), .B0(n65), .Y(n70) );
  OA21X2 U14 ( .A0(n44), .A1(n45), .B0(n41), .Y(n46) );
  OA21X2 U15 ( .A0(n20), .A1(n21), .B0(n17), .Y(n22) );
  OAI21X2 U16 ( .A0(n124), .A1(n122), .B0(n121), .Y(n130) );
  OA21X2 U17 ( .A0(n116), .A1(n117), .B0(n113), .Y(n118) );
  MXI2XL U18 ( .A(n120), .B(n119), .S0(n118), .Y(n121) );
  MXI2XL U19 ( .A(n8), .B(n7), .S0(n6), .Y(n9) );
  MXI2XL U20 ( .A(n16), .B(n15), .S0(n14), .Y(n17) );
  MXI2XL U21 ( .A(n24), .B(n23), .S0(n22), .Y(n25) );
  MXI2XL U22 ( .A(n32), .B(n31), .S0(n30), .Y(n33) );
  MXI2XL U23 ( .A(n40), .B(n39), .S0(n38), .Y(n41) );
  MXI2XL U24 ( .A(n48), .B(n47), .S0(n46), .Y(n49) );
  MXI2XL U25 ( .A(n56), .B(n55), .S0(n54), .Y(n57) );
  MXI2XL U26 ( .A(n64), .B(n63), .S0(n62), .Y(n65) );
  MXI2XL U27 ( .A(n72), .B(n71), .S0(n70), .Y(n73) );
  MXI2XL U28 ( .A(n80), .B(n79), .S0(n78), .Y(n81) );
  MXI2XL U29 ( .A(n88), .B(n87), .S0(n86), .Y(n89) );
  MXI2XL U30 ( .A(n96), .B(n95), .S0(n94), .Y(n97) );
  MXI2XL U31 ( .A(n104), .B(n103), .S0(n102), .Y(n105) );
  MXI2XL U32 ( .A(n112), .B(n111), .S0(n110), .Y(n113) );
  XNOR2XL U33 ( .A(n122), .B(n124), .Y(n123) );
  CLKINVX1 U34 ( .A(\u_div/SumTmp[17][0] ), .Y(n128) );
  NAND2X1 U35 ( .A(n129), .B(\u_div/SumTmp[19][0] ), .Y(n1) );
  CLKMX2X2 U36 ( .A(n128), .B(\u_div/SumTmp[17][0] ), .S0(n1), .Y(n2) );
  XOR2X1 U37 ( .A(\u_div/SumTmp[16][0] ), .B(n2), .Y(n3) );
  MXI2X1 U38 ( .A(\u_div/SumTmp[16][2] ), .B(\u_div/SumTmp[18][0] ), .S0(n1), 
        .Y(n4) );
  NAND2X1 U39 ( .A(\u_div/SumTmp[16][0] ), .B(n2), .Y(n5) );
  MXI2X1 U40 ( .A(n3), .B(n2), .S0(n6), .Y(n12) );
  XNOR2X1 U41 ( .A(\u_div/SumTmp[16][0] ), .B(n6), .Y(n10) );
  NAND2X1 U42 ( .A(\u_div/SumTmp[15][0] ), .B(n10), .Y(n13) );
  CLKINVX1 U43 ( .A(n4), .Y(n7) );
  XNOR2X1 U44 ( .A(n5), .B(n7), .Y(n8) );
  XNOR2X1 U45 ( .A(\u_div/SumTmp[15][0] ), .B(n14), .Y(n18) );
  XOR2X1 U46 ( .A(n18), .B(\u_div/SumTmp[14][0] ), .Y(n19) );
  XOR2X1 U47 ( .A(n10), .B(\u_div/SumTmp[15][0] ), .Y(n11) );
  MXI2X1 U48 ( .A(n11), .B(n10), .S0(n14), .Y(n20) );
  NAND2X1 U49 ( .A(\u_div/SumTmp[14][0] ), .B(n18), .Y(n21) );
  CLKINVX1 U50 ( .A(n12), .Y(n15) );
  XNOR2X1 U51 ( .A(n13), .B(n15), .Y(n16) );
  MXI2X1 U52 ( .A(n19), .B(n18), .S0(n22), .Y(n28) );
  XNOR2X1 U53 ( .A(\u_div/SumTmp[14][0] ), .B(n22), .Y(n26) );
  NAND2X1 U54 ( .A(\u_div/SumTmp[13][0] ), .B(n26), .Y(n29) );
  CLKINVX1 U55 ( .A(n20), .Y(n23) );
  XNOR2X1 U56 ( .A(n21), .B(n23), .Y(n24) );
  XNOR2X1 U57 ( .A(\u_div/SumTmp[13][0] ), .B(n30), .Y(n34) );
  XOR2X1 U58 ( .A(n34), .B(\u_div/SumTmp[12][0] ), .Y(n35) );
  XOR2X1 U59 ( .A(n26), .B(\u_div/SumTmp[13][0] ), .Y(n27) );
  MXI2X1 U60 ( .A(n27), .B(n26), .S0(n30), .Y(n36) );
  NAND2X1 U61 ( .A(\u_div/SumTmp[12][0] ), .B(n34), .Y(n37) );
  CLKINVX1 U62 ( .A(n28), .Y(n31) );
  XNOR2X1 U63 ( .A(n29), .B(n31), .Y(n32) );
  MXI2X1 U64 ( .A(n35), .B(n34), .S0(n38), .Y(n44) );
  XNOR2X1 U65 ( .A(\u_div/SumTmp[12][0] ), .B(n38), .Y(n42) );
  NAND2X1 U66 ( .A(\u_div/SumTmp[11][0] ), .B(n42), .Y(n45) );
  CLKINVX1 U67 ( .A(n36), .Y(n39) );
  XNOR2X1 U68 ( .A(n37), .B(n39), .Y(n40) );
  XNOR2X1 U69 ( .A(\u_div/SumTmp[11][0] ), .B(n46), .Y(n50) );
  XOR2X1 U70 ( .A(n50), .B(\u_div/SumTmp[10][0] ), .Y(n51) );
  XOR2X1 U71 ( .A(n42), .B(\u_div/SumTmp[11][0] ), .Y(n43) );
  MXI2X1 U72 ( .A(n43), .B(n42), .S0(n46), .Y(n52) );
  NAND2X1 U73 ( .A(\u_div/SumTmp[10][0] ), .B(n50), .Y(n53) );
  CLKINVX1 U74 ( .A(n44), .Y(n47) );
  XNOR2X1 U75 ( .A(n45), .B(n47), .Y(n48) );
  MXI2X1 U76 ( .A(n51), .B(n50), .S0(n54), .Y(n60) );
  XNOR2X1 U77 ( .A(\u_div/SumTmp[10][0] ), .B(n54), .Y(n58) );
  NAND2X1 U78 ( .A(\u_div/SumTmp[9][0] ), .B(n58), .Y(n61) );
  CLKINVX1 U79 ( .A(n52), .Y(n55) );
  XNOR2X1 U80 ( .A(n53), .B(n55), .Y(n56) );
  XNOR2X1 U81 ( .A(\u_div/SumTmp[9][0] ), .B(n62), .Y(n66) );
  XOR2X1 U82 ( .A(n66), .B(\u_div/SumTmp[8][0] ), .Y(n67) );
  XOR2X1 U83 ( .A(n58), .B(\u_div/SumTmp[9][0] ), .Y(n59) );
  MXI2X1 U84 ( .A(n59), .B(n58), .S0(n62), .Y(n68) );
  NAND2X1 U85 ( .A(\u_div/SumTmp[8][0] ), .B(n66), .Y(n69) );
  CLKINVX1 U86 ( .A(n60), .Y(n63) );
  XNOR2X1 U87 ( .A(n61), .B(n63), .Y(n64) );
  MXI2X1 U88 ( .A(n67), .B(n66), .S0(n70), .Y(n76) );
  XNOR2X1 U89 ( .A(\u_div/SumTmp[8][0] ), .B(n70), .Y(n74) );
  NAND2X1 U90 ( .A(\u_div/SumTmp[7][0] ), .B(n74), .Y(n77) );
  CLKINVX1 U91 ( .A(n68), .Y(n71) );
  XNOR2X1 U92 ( .A(n69), .B(n71), .Y(n72) );
  XNOR2X1 U93 ( .A(\u_div/SumTmp[7][0] ), .B(n78), .Y(n82) );
  XOR2X1 U94 ( .A(n82), .B(\u_div/SumTmp[6][0] ), .Y(n83) );
  XOR2X1 U95 ( .A(n74), .B(\u_div/SumTmp[7][0] ), .Y(n75) );
  MXI2X1 U96 ( .A(n75), .B(n74), .S0(n78), .Y(n84) );
  NAND2X1 U97 ( .A(\u_div/SumTmp[6][0] ), .B(n82), .Y(n85) );
  CLKINVX1 U98 ( .A(n76), .Y(n79) );
  XNOR2X1 U99 ( .A(n77), .B(n79), .Y(n80) );
  MXI2X1 U100 ( .A(n83), .B(n82), .S0(n86), .Y(n92) );
  XNOR2X1 U101 ( .A(\u_div/SumTmp[6][0] ), .B(n86), .Y(n90) );
  NAND2X1 U102 ( .A(\u_div/SumTmp[5][0] ), .B(n90), .Y(n93) );
  CLKINVX1 U103 ( .A(n84), .Y(n87) );
  XNOR2X1 U104 ( .A(n85), .B(n87), .Y(n88) );
  XNOR2X1 U105 ( .A(\u_div/SumTmp[5][0] ), .B(n94), .Y(n98) );
  XOR2X1 U106 ( .A(n98), .B(\u_div/SumTmp[4][0] ), .Y(n99) );
  XOR2X1 U107 ( .A(n90), .B(\u_div/SumTmp[5][0] ), .Y(n91) );
  MXI2X1 U108 ( .A(n91), .B(n90), .S0(n94), .Y(n100) );
  NAND2X1 U109 ( .A(\u_div/SumTmp[4][0] ), .B(n98), .Y(n101) );
  CLKINVX1 U110 ( .A(n92), .Y(n95) );
  XNOR2X1 U111 ( .A(n93), .B(n95), .Y(n96) );
  MXI2X1 U112 ( .A(n99), .B(n98), .S0(n102), .Y(n108) );
  XNOR2X1 U113 ( .A(\u_div/SumTmp[4][0] ), .B(n102), .Y(n106) );
  NAND2X1 U114 ( .A(\u_div/SumTmp[3][0] ), .B(n106), .Y(n109) );
  CLKINVX1 U115 ( .A(n100), .Y(n103) );
  XNOR2X1 U116 ( .A(n101), .B(n103), .Y(n104) );
  XNOR2X1 U117 ( .A(\u_div/SumTmp[3][0] ), .B(n110), .Y(n114) );
  XOR2X1 U118 ( .A(n114), .B(\u_div/SumTmp[2][0] ), .Y(n115) );
  XOR2X1 U119 ( .A(n106), .B(\u_div/SumTmp[3][0] ), .Y(n107) );
  MXI2X1 U120 ( .A(n107), .B(n106), .S0(n110), .Y(n116) );
  NAND2X1 U121 ( .A(\u_div/SumTmp[2][0] ), .B(n114), .Y(n117) );
  CLKINVX1 U122 ( .A(n108), .Y(n111) );
  XNOR2X1 U123 ( .A(n109), .B(n111), .Y(n112) );
  XOR2X1 U124 ( .A(\u_div/SumTmp[2][0] ), .B(n118), .Y(n127) );
  NAND2BX1 U125 ( .AN(n127), .B(\u_div/SumTmp[1][0] ), .Y(n122) );
  CLKINVX1 U126 ( .A(n116), .Y(n119) );
  XNOR2X1 U127 ( .A(n117), .B(n119), .Y(n120) );
  CLKINVX1 U128 ( .A(\u_div/SumTmp[1][0] ), .Y(n125) );
  XNOR2X1 U129 ( .A(n125), .B(n130), .Y(remainder[1]) );
  MXI2X1 U130 ( .A(n124), .B(n123), .S0(n130), .Y(remainder[3]) );
  XNOR2X1 U131 ( .A(n125), .B(n127), .Y(n126) );
  MXI2X1 U132 ( .A(n127), .B(n126), .S0(n130), .Y(remainder[2]) );
  NOR2BX1 U133 ( .AN(\u_div/SumTmp[18][0] ), .B(n128), .Y(n129) );
  XOR2X1 U134 ( .A(\u_div/SumTmp[18][0] ), .B(\u_div/SumTmp[17][0] ), .Y(
        \u_div/SumTmp[16][2] ) );
endmodule


module CONT_DW_div_uns_59 ( a, b, quotient, remainder, divide_by_0 );
  input [8:0] a;
  input [4:0] b;
  output [8:0] quotient;
  output [4:0] remainder;
  output divide_by_0;
  wire   n31, n32, n33, n34, \u_div/SumTmp[0][0] , \u_div/SumTmp[1][0] ,
         \u_div/SumTmp[2][0] , \u_div/SumTmp[3][0] , \u_div/SumTmp[4][0] ,
         \u_div/CryTmp[0][4] , \u_div/CryTmp[1][4] , \u_div/CryTmp[2][4] ,
         \u_div/CryTmp[3][4] , \u_div/CryTmp[4][4] , \u_div/PartRem[1][4] ,
         \u_div/PartRem[1][5] , \u_div/PartRem[2][4] , \u_div/PartRem[2][5] ,
         \u_div/PartRem[3][4] , \u_div/PartRem[3][5] , \u_div/PartRem[4][4] ,
         \u_div/PartRem[4][5] , \u_div/PartRem[5][4] , \u_div/PartRem[7][1] ,
         \u_div/PartRem[8][1] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30;
  assign \u_div/SumTmp[0][0]  = a[0];
  assign \u_div/SumTmp[1][0]  = a[1];
  assign \u_div/SumTmp[2][0]  = a[2];
  assign \u_div/SumTmp[3][0]  = a[3];
  assign \u_div/SumTmp[4][0]  = a[4];
  assign \u_div/PartRem[7][1]  = a[7];
  assign \u_div/PartRem[8][1]  = a[8];

  CLKMX2X2 U1 ( .A(a[5]), .B(a[5]), .S0(n13), .Y(n1) );
  CLKMX2X2 U2 ( .A(n5), .B(n5), .S0(n32), .Y(n2) );
  CLKMX2X2 U3 ( .A(n17), .B(n17), .S0(n31), .Y(n3) );
  XNOR2X1 U4 ( .A(\u_div/PartRem[1][4] ), .B(\u_div/CryTmp[0][4] ), .Y(n4) );
  CLKMX2X2 U5 ( .A(\u_div/SumTmp[3][0] ), .B(\u_div/SumTmp[3][0] ), .S0(n31), 
        .Y(n5) );
  OR2X2 U6 ( .A(\u_div/PartRem[2][5] ), .B(n8), .Y(n33) );
  OR2X2 U7 ( .A(\u_div/PartRem[1][5] ), .B(n6), .Y(n34) );
  CLKBUFX3 U8 ( .A(n19), .Y(remainder[3]) );
  OR2X2 U9 ( .A(\u_div/PartRem[3][5] ), .B(n7), .Y(n32) );
  OR2X2 U10 ( .A(\u_div/PartRem[4][5] ), .B(n9), .Y(n31) );
  MXI2X1 U11 ( .A(n24), .B(n10), .S0(n32), .Y(\u_div/PartRem[2][5] ) );
  MXI2X1 U12 ( .A(n26), .B(n11), .S0(n33), .Y(\u_div/PartRem[1][5] ) );
  CLKINVX1 U13 ( .A(n24), .Y(\u_div/PartRem[3][4] ) );
  CLKINVX1 U14 ( .A(n26), .Y(\u_div/PartRem[2][4] ) );
  CLKINVX1 U15 ( .A(n28), .Y(\u_div/PartRem[1][4] ) );
  AND2X2 U16 ( .A(\u_div/CryTmp[0][4] ), .B(\u_div/PartRem[1][4] ), .Y(n6) );
  CLKBUFX3 U17 ( .A(n20), .Y(remainder[4]) );
  MXI2X1 U18 ( .A(n28), .B(n4), .S0(n34), .Y(n20) );
  MXI2X1 U19 ( .A(n22), .B(n12), .S0(n31), .Y(\u_div/PartRem[3][5] ) );
  CLKMX2X2 U20 ( .A(n25), .B(\u_div/CryTmp[3][4] ), .S0(n31), .Y(n24) );
  CLKMX2X2 U21 ( .A(n27), .B(\u_div/CryTmp[2][4] ), .S0(n32), .Y(n26) );
  CLKMX2X2 U22 ( .A(n30), .B(\u_div/CryTmp[1][4] ), .S0(n33), .Y(n28) );
  CLKINVX1 U23 ( .A(n29), .Y(\u_div/CryTmp[0][4] ) );
  CLKINVX1 U24 ( .A(n22), .Y(\u_div/PartRem[4][4] ) );
  AND2X2 U25 ( .A(\u_div/CryTmp[2][4] ), .B(\u_div/PartRem[3][4] ), .Y(n7) );
  AND2X2 U26 ( .A(\u_div/CryTmp[1][4] ), .B(\u_div/PartRem[2][4] ), .Y(n8) );
  AND2X2 U27 ( .A(\u_div/CryTmp[3][4] ), .B(\u_div/PartRem[4][4] ), .Y(n9) );
  XNOR2X1 U28 ( .A(\u_div/PartRem[3][4] ), .B(\u_div/CryTmp[2][4] ), .Y(n10)
         );
  XNOR2X1 U29 ( .A(\u_div/PartRem[2][4] ), .B(\u_div/CryTmp[1][4] ), .Y(n11)
         );
  XNOR2X1 U30 ( .A(\u_div/PartRem[4][4] ), .B(\u_div/CryTmp[3][4] ), .Y(n12)
         );
  MXI2X1 U31 ( .A(n21), .B(n14), .S0(n13), .Y(\u_div/PartRem[4][5] ) );
  CLKMX2X2 U32 ( .A(n23), .B(\u_div/CryTmp[4][4] ), .S0(n13), .Y(n22) );
  MXI2X1 U33 ( .A(n2), .B(n2), .S0(n33), .Y(n29) );
  CLKINVX1 U34 ( .A(n25), .Y(\u_div/CryTmp[3][4] ) );
  MXI2X1 U35 ( .A(a[6]), .B(a[6]), .S0(n13), .Y(n25) );
  CLKINVX1 U36 ( .A(n27), .Y(\u_div/CryTmp[2][4] ) );
  MXI2X1 U37 ( .A(n1), .B(n1), .S0(n31), .Y(n27) );
  CLKINVX1 U38 ( .A(n30), .Y(\u_div/CryTmp[1][4] ) );
  MXI2X1 U39 ( .A(n3), .B(n3), .S0(n32), .Y(n30) );
  AND2X2 U40 ( .A(\u_div/CryTmp[4][4] ), .B(\u_div/PartRem[5][4] ), .Y(n13) );
  CLKINVX1 U41 ( .A(n21), .Y(\u_div/PartRem[5][4] ) );
  XNOR2X1 U42 ( .A(\u_div/PartRem[5][4] ), .B(\u_div/CryTmp[4][4] ), .Y(n14)
         );
  CLKMX2X2 U43 ( .A(n15), .B(n15), .S0(n34), .Y(remainder[2]) );
  CLKMX2X2 U44 ( .A(n18), .B(n18), .S0(n33), .Y(n15) );
  CLKINVX1 U45 ( .A(\u_div/PartRem[8][1] ), .Y(n21) );
  CLKINVX1 U46 ( .A(n23), .Y(\u_div/CryTmp[4][4] ) );
  CLKINVX1 U47 ( .A(\u_div/PartRem[7][1] ), .Y(n23) );
  CLKMX2X2 U48 ( .A(\u_div/SumTmp[0][0] ), .B(\u_div/SumTmp[0][0] ), .S0(n34), 
        .Y(remainder[0]) );
  CLKMX2X2 U49 ( .A(n16), .B(n16), .S0(n34), .Y(remainder[1]) );
  CLKMX2X2 U50 ( .A(\u_div/SumTmp[1][0] ), .B(\u_div/SumTmp[1][0] ), .S0(n33), 
        .Y(n16) );
  CLKMX2X2 U51 ( .A(\u_div/SumTmp[4][0] ), .B(\u_div/SumTmp[4][0] ), .S0(n13), 
        .Y(n17) );
  CLKMX2X2 U52 ( .A(\u_div/SumTmp[2][0] ), .B(\u_div/SumTmp[2][0] ), .S0(n32), 
        .Y(n18) );
  MXI2X1 U53 ( .A(n29), .B(\u_div/CryTmp[0][4] ), .S0(n34), .Y(n19) );
endmodule


module CONT_DW_div_uns_71 ( a, b, quotient, remainder, divide_by_0 );
  input [19:0] a;
  input [4:0] b;
  output [19:0] quotient;
  output [4:0] remainder;
  output divide_by_0;
  wire   n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         \u_div/SumTmp[0][0] , \u_div/SumTmp[1][0] , \u_div/SumTmp[2][0] ,
         \u_div/SumTmp[3][0] , \u_div/SumTmp[4][0] , \u_div/SumTmp[5][0] ,
         \u_div/SumTmp[6][0] , \u_div/SumTmp[7][0] , \u_div/SumTmp[8][0] ,
         \u_div/SumTmp[9][0] , \u_div/SumTmp[10][0] , \u_div/SumTmp[11][0] ,
         \u_div/SumTmp[12][0] , \u_div/CryTmp[0][4] , \u_div/CryTmp[1][4] ,
         \u_div/CryTmp[2][4] , \u_div/CryTmp[3][4] , \u_div/CryTmp[4][4] ,
         \u_div/CryTmp[5][4] , \u_div/CryTmp[6][4] , \u_div/CryTmp[7][4] ,
         \u_div/CryTmp[8][4] , \u_div/CryTmp[9][4] , \u_div/CryTmp[10][4] ,
         \u_div/CryTmp[11][4] , \u_div/PartRem[1][4] , \u_div/PartRem[1][5] ,
         \u_div/PartRem[2][4] , \u_div/PartRem[2][5] , \u_div/PartRem[3][4] ,
         \u_div/PartRem[3][5] , \u_div/PartRem[4][4] , \u_div/PartRem[4][5] ,
         \u_div/PartRem[5][4] , \u_div/PartRem[5][5] , \u_div/PartRem[6][4] ,
         \u_div/PartRem[6][5] , \u_div/PartRem[7][4] , \u_div/PartRem[7][5] ,
         \u_div/PartRem[8][4] , \u_div/PartRem[8][5] , \u_div/PartRem[9][4] ,
         \u_div/PartRem[9][5] , \u_div/PartRem[10][4] , \u_div/PartRem[10][5] ,
         \u_div/PartRem[11][4] , \u_div/PartRem[11][5] ,
         \u_div/PartRem[12][4] , \u_div/PartRem[12][5] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77;
  assign \u_div/SumTmp[0][0]  = a[0];
  assign \u_div/SumTmp[1][0]  = a[1];
  assign \u_div/SumTmp[2][0]  = a[2];
  assign \u_div/SumTmp[3][0]  = a[3];
  assign \u_div/SumTmp[4][0]  = a[4];
  assign \u_div/SumTmp[5][0]  = a[5];
  assign \u_div/SumTmp[6][0]  = a[6];
  assign \u_div/SumTmp[7][0]  = a[7];
  assign \u_div/SumTmp[8][0]  = a[8];
  assign \u_div/SumTmp[9][0]  = a[9];
  assign \u_div/SumTmp[10][0]  = a[10];
  assign \u_div/SumTmp[11][0]  = a[11];
  assign \u_div/SumTmp[12][0]  = a[12];

  CLKMX2X2 U1 ( .A(n35), .B(n35), .S0(n86), .Y(n1) );
  CLKMX2X2 U2 ( .A(n36), .B(n36), .S0(n85), .Y(n2) );
  CLKMX2X2 U3 ( .A(n37), .B(n37), .S0(n84), .Y(n3) );
  CLKMX2X2 U4 ( .A(n38), .B(n38), .S0(n83), .Y(n4) );
  CLKMX2X2 U5 ( .A(n39), .B(n39), .S0(n82), .Y(n5) );
  CLKMX2X2 U6 ( .A(n40), .B(n40), .S0(n81), .Y(n6) );
  CLKMX2X2 U7 ( .A(n41), .B(n41), .S0(n80), .Y(n7) );
  CLKMX2X2 U8 ( .A(n42), .B(n42), .S0(n79), .Y(n8) );
  CLKMX2X2 U9 ( .A(n43), .B(n43), .S0(n78), .Y(n9) );
  CLKMX2X2 U10 ( .A(a[13]), .B(a[13]), .S0(n44), .Y(n10) );
  XNOR2X1 U11 ( .A(\u_div/PartRem[1][4] ), .B(\u_div/CryTmp[0][4] ), .Y(n11)
         );
  MX2XL U12 ( .A(\u_div/SumTmp[4][0] ), .B(\u_div/SumTmp[4][0] ), .S0(n85), 
        .Y(n35) );
  MX2XL U13 ( .A(\u_div/SumTmp[5][0] ), .B(\u_div/SumTmp[5][0] ), .S0(n84), 
        .Y(n36) );
  MX2XL U14 ( .A(\u_div/SumTmp[6][0] ), .B(\u_div/SumTmp[6][0] ), .S0(n83), 
        .Y(n37) );
  MX2XL U15 ( .A(\u_div/SumTmp[7][0] ), .B(\u_div/SumTmp[7][0] ), .S0(n82), 
        .Y(n38) );
  MX2XL U16 ( .A(\u_div/SumTmp[8][0] ), .B(\u_div/SumTmp[8][0] ), .S0(n81), 
        .Y(n39) );
  MX2XL U17 ( .A(\u_div/SumTmp[9][0] ), .B(\u_div/SumTmp[9][0] ), .S0(n80), 
        .Y(n40) );
  MX2XL U18 ( .A(\u_div/SumTmp[10][0] ), .B(\u_div/SumTmp[10][0] ), .S0(n79), 
        .Y(n41) );
  MX2XL U19 ( .A(\u_div/SumTmp[11][0] ), .B(\u_div/SumTmp[11][0] ), .S0(n78), 
        .Y(n42) );
  MX2XL U20 ( .A(\u_div/SumTmp[12][0] ), .B(\u_div/SumTmp[12][0] ), .S0(n44), 
        .Y(n43) );
  OR2X2 U21 ( .A(\u_div/PartRem[1][5] ), .B(n12), .Y(n89) );
  OR2X2 U22 ( .A(\u_div/PartRem[2][5] ), .B(n13), .Y(n88) );
  OR2X2 U23 ( .A(\u_div/PartRem[3][5] ), .B(n14), .Y(n87) );
  OR2X2 U24 ( .A(\u_div/PartRem[4][5] ), .B(n18), .Y(n86) );
  OR2X2 U25 ( .A(\u_div/PartRem[5][5] ), .B(n19), .Y(n85) );
  OR2X2 U26 ( .A(\u_div/PartRem[6][5] ), .B(n22), .Y(n84) );
  OR2X2 U27 ( .A(\u_div/PartRem[7][5] ), .B(n23), .Y(n83) );
  OR2X2 U28 ( .A(\u_div/PartRem[8][5] ), .B(n26), .Y(n82) );
  OR2X2 U29 ( .A(\u_div/PartRem[9][5] ), .B(n27), .Y(n81) );
  OR2X2 U30 ( .A(\u_div/PartRem[10][5] ), .B(n30), .Y(n80) );
  OR2X2 U31 ( .A(\u_div/PartRem[11][5] ), .B(n31), .Y(n79) );
  OR2X2 U32 ( .A(\u_div/PartRem[12][5] ), .B(n34), .Y(n78) );
  MXI2X1 U33 ( .A(n60), .B(n15), .S0(n88), .Y(\u_div/PartRem[1][5] ) );
  AND2X2 U34 ( .A(\u_div/CryTmp[0][4] ), .B(\u_div/PartRem[1][4] ), .Y(n12) );
  MXI2X1 U35 ( .A(n58), .B(n16), .S0(n87), .Y(\u_div/PartRem[2][5] ) );
  CLKINVX1 U36 ( .A(n62), .Y(\u_div/PartRem[1][4] ) );
  MXI2X1 U37 ( .A(n56), .B(n17), .S0(n86), .Y(\u_div/PartRem[3][5] ) );
  CLKINVX1 U38 ( .A(n60), .Y(\u_div/PartRem[2][4] ) );
  MXI2X1 U39 ( .A(n54), .B(n20), .S0(n85), .Y(\u_div/PartRem[4][5] ) );
  CLKINVX1 U40 ( .A(n58), .Y(\u_div/PartRem[3][4] ) );
  MXI2X1 U41 ( .A(n52), .B(n21), .S0(n84), .Y(\u_div/PartRem[5][5] ) );
  CLKINVX1 U42 ( .A(n56), .Y(\u_div/PartRem[4][4] ) );
  MXI2X1 U43 ( .A(n50), .B(n24), .S0(n83), .Y(\u_div/PartRem[6][5] ) );
  CLKINVX1 U44 ( .A(n54), .Y(\u_div/PartRem[5][4] ) );
  MXI2X1 U45 ( .A(n48), .B(n25), .S0(n82), .Y(\u_div/PartRem[7][5] ) );
  CLKINVX1 U46 ( .A(n52), .Y(\u_div/PartRem[6][4] ) );
  MXI2X1 U47 ( .A(n47), .B(n28), .S0(n81), .Y(\u_div/PartRem[8][5] ) );
  CLKINVX1 U48 ( .A(n50), .Y(\u_div/PartRem[7][4] ) );
  MXI2X1 U49 ( .A(n46), .B(n29), .S0(n80), .Y(\u_div/PartRem[9][5] ) );
  CLKINVX1 U50 ( .A(n48), .Y(\u_div/PartRem[8][4] ) );
  CLKINVX1 U51 ( .A(n47), .Y(\u_div/PartRem[9][4] ) );
  CLKINVX1 U52 ( .A(n46), .Y(\u_div/PartRem[10][4] ) );
  CLKINVX1 U53 ( .A(n63), .Y(\u_div/CryTmp[0][4] ) );
  MXI2X1 U54 ( .A(\u_div/CryTmp[1][4] ), .B(n73), .S0(n88), .Y(n62) );
  AND2X2 U55 ( .A(\u_div/CryTmp[1][4] ), .B(\u_div/PartRem[2][4] ), .Y(n13) );
  CLKMX2X2 U56 ( .A(n61), .B(\u_div/CryTmp[2][4] ), .S0(n87), .Y(n60) );
  AND2X2 U57 ( .A(\u_div/CryTmp[2][4] ), .B(\u_div/PartRem[3][4] ), .Y(n14) );
  XNOR2X1 U58 ( .A(\u_div/PartRem[2][4] ), .B(\u_div/CryTmp[1][4] ), .Y(n15)
         );
  XNOR2X1 U59 ( .A(\u_div/PartRem[3][4] ), .B(\u_div/CryTmp[2][4] ), .Y(n16)
         );
  CLKMX2X2 U60 ( .A(n59), .B(\u_div/CryTmp[3][4] ), .S0(n86), .Y(n58) );
  XNOR2X1 U61 ( .A(\u_div/PartRem[4][4] ), .B(\u_div/CryTmp[3][4] ), .Y(n17)
         );
  AND2X2 U62 ( .A(\u_div/CryTmp[3][4] ), .B(\u_div/PartRem[4][4] ), .Y(n18) );
  CLKMX2X2 U63 ( .A(n57), .B(\u_div/CryTmp[4][4] ), .S0(n85), .Y(n56) );
  AND2X2 U64 ( .A(\u_div/CryTmp[4][4] ), .B(\u_div/PartRem[5][4] ), .Y(n19) );
  XNOR2X1 U65 ( .A(\u_div/PartRem[5][4] ), .B(\u_div/CryTmp[4][4] ), .Y(n20)
         );
  CLKMX2X2 U66 ( .A(n55), .B(\u_div/CryTmp[5][4] ), .S0(n84), .Y(n54) );
  XNOR2X1 U67 ( .A(\u_div/PartRem[6][4] ), .B(\u_div/CryTmp[5][4] ), .Y(n21)
         );
  AND2X2 U68 ( .A(\u_div/CryTmp[5][4] ), .B(\u_div/PartRem[6][4] ), .Y(n22) );
  CLKMX2X2 U69 ( .A(n53), .B(\u_div/CryTmp[6][4] ), .S0(n83), .Y(n52) );
  AND2X2 U70 ( .A(\u_div/CryTmp[6][4] ), .B(\u_div/PartRem[7][4] ), .Y(n23) );
  XNOR2X1 U71 ( .A(\u_div/PartRem[7][4] ), .B(\u_div/CryTmp[6][4] ), .Y(n24)
         );
  CLKMX2X2 U72 ( .A(n51), .B(\u_div/CryTmp[7][4] ), .S0(n82), .Y(n50) );
  XNOR2X1 U73 ( .A(\u_div/PartRem[8][4] ), .B(\u_div/CryTmp[7][4] ), .Y(n25)
         );
  AND2X2 U74 ( .A(\u_div/CryTmp[7][4] ), .B(\u_div/PartRem[8][4] ), .Y(n26) );
  CLKMX2X2 U75 ( .A(n49), .B(\u_div/CryTmp[8][4] ), .S0(n81), .Y(n48) );
  AND2X2 U76 ( .A(\u_div/CryTmp[8][4] ), .B(\u_div/PartRem[9][4] ), .Y(n27) );
  XNOR2X1 U77 ( .A(\u_div/PartRem[9][4] ), .B(\u_div/CryTmp[8][4] ), .Y(n28)
         );
  MXI2X1 U78 ( .A(n69), .B(n32), .S0(n79), .Y(\u_div/PartRem[10][5] ) );
  CLKMX2X2 U79 ( .A(n72), .B(\u_div/CryTmp[9][4] ), .S0(n80), .Y(n47) );
  XNOR2X1 U80 ( .A(\u_div/PartRem[10][4] ), .B(\u_div/CryTmp[9][4] ), .Y(n29)
         );
  AND2X2 U81 ( .A(\u_div/CryTmp[9][4] ), .B(\u_div/PartRem[10][4] ), .Y(n30)
         );
  CLKMX2X2 U82 ( .A(n71), .B(\u_div/CryTmp[10][4] ), .S0(n79), .Y(n46) );
  AND2X2 U83 ( .A(\u_div/CryTmp[10][4] ), .B(\u_div/PartRem[11][4] ), .Y(n31)
         );
  XNOR2X1 U84 ( .A(\u_div/PartRem[11][4] ), .B(\u_div/CryTmp[10][4] ), .Y(n32)
         );
  CLKINVX1 U85 ( .A(n69), .Y(\u_div/PartRem[11][4] ) );
  MXI2X1 U86 ( .A(n64), .B(n64), .S0(n89), .Y(remainder[2]) );
  MXI2X1 U87 ( .A(n63), .B(\u_div/CryTmp[0][4] ), .S0(n89), .Y(remainder[3])
         );
  MXI2X1 U88 ( .A(n62), .B(n11), .S0(n89), .Y(remainder[4]) );
  CLKMX2X2 U89 ( .A(n74), .B(n74), .S0(n88), .Y(n63) );
  CLKMX2X2 U90 ( .A(n75), .B(n75), .S0(n87), .Y(n74) );
  CLKINVX1 U91 ( .A(n73), .Y(\u_div/CryTmp[1][4] ) );
  MXI2X1 U92 ( .A(n1), .B(n1), .S0(n87), .Y(n73) );
  CLKINVX1 U93 ( .A(n61), .Y(\u_div/CryTmp[2][4] ) );
  MXI2X1 U94 ( .A(n2), .B(n2), .S0(n86), .Y(n61) );
  CLKINVX1 U95 ( .A(n59), .Y(\u_div/CryTmp[3][4] ) );
  MXI2X1 U96 ( .A(n3), .B(n3), .S0(n85), .Y(n59) );
  CLKINVX1 U97 ( .A(n57), .Y(\u_div/CryTmp[4][4] ) );
  MXI2X1 U98 ( .A(n4), .B(n4), .S0(n84), .Y(n57) );
  CLKINVX1 U99 ( .A(n55), .Y(\u_div/CryTmp[5][4] ) );
  MXI2X1 U100 ( .A(n5), .B(n5), .S0(n83), .Y(n55) );
  CLKINVX1 U101 ( .A(n53), .Y(\u_div/CryTmp[6][4] ) );
  MXI2X1 U102 ( .A(n6), .B(n6), .S0(n82), .Y(n53) );
  CLKINVX1 U103 ( .A(n51), .Y(\u_div/CryTmp[7][4] ) );
  MXI2X1 U104 ( .A(n7), .B(n7), .S0(n81), .Y(n51) );
  CLKINVX1 U105 ( .A(n49), .Y(\u_div/CryTmp[8][4] ) );
  MXI2X1 U106 ( .A(n8), .B(n8), .S0(n80), .Y(n49) );
  CLKINVX1 U107 ( .A(n72), .Y(\u_div/CryTmp[9][4] ) );
  MXI2X1 U108 ( .A(n9), .B(n9), .S0(n79), .Y(n72) );
  MXI2X1 U109 ( .A(n67), .B(n33), .S0(n78), .Y(\u_div/PartRem[11][5] ) );
  CLKINVX1 U110 ( .A(n71), .Y(\u_div/CryTmp[10][4] ) );
  MXI2X1 U111 ( .A(n10), .B(n10), .S0(n78), .Y(n71) );
  CLKMX2X2 U112 ( .A(n70), .B(\u_div/CryTmp[11][4] ), .S0(n78), .Y(n69) );
  XNOR2X1 U113 ( .A(\u_div/PartRem[12][4] ), .B(\u_div/CryTmp[11][4] ), .Y(n33) );
  AND2X2 U114 ( .A(\u_div/CryTmp[11][4] ), .B(\u_div/PartRem[12][4] ), .Y(n34)
         );
  CLKINVX1 U115 ( .A(n67), .Y(\u_div/PartRem[12][4] ) );
  MXI2XL U116 ( .A(n65), .B(n65), .S0(n89), .Y(remainder[1]) );
  MXI2X1 U117 ( .A(\u_div/SumTmp[1][0] ), .B(\u_div/SumTmp[1][0] ), .S0(n88), 
        .Y(n65) );
  CLKMX2X2 U118 ( .A(n76), .B(n76), .S0(n88), .Y(n64) );
  MXI2X1 U119 ( .A(\u_div/SumTmp[2][0] ), .B(\u_div/SumTmp[2][0] ), .S0(n87), 
        .Y(n76) );
  MXI2X1 U120 ( .A(\u_div/SumTmp[3][0] ), .B(\u_div/SumTmp[3][0] ), .S0(n86), 
        .Y(n75) );
  MXI2X1 U121 ( .A(n66), .B(n45), .S0(n44), .Y(\u_div/PartRem[12][5] ) );
  CLKINVX1 U122 ( .A(n70), .Y(\u_div/CryTmp[11][4] ) );
  MXI2X1 U123 ( .A(a[14]), .B(a[14]), .S0(n44), .Y(n70) );
  CLKMX2X2 U124 ( .A(n68), .B(a[15]), .S0(n44), .Y(n67) );
  AND2X2 U125 ( .A(a[15]), .B(a[16]), .Y(n44) );
  XNOR2X1 U126 ( .A(a[16]), .B(a[15]), .Y(n45) );
  MXI2X1 U127 ( .A(n77), .B(n77), .S0(n89), .Y(remainder[0]) );
  CLKINVX1 U128 ( .A(\u_div/SumTmp[0][0] ), .Y(n77) );
  INVXL U129 ( .A(a[15]), .Y(n68) );
  INVXL U130 ( .A(a[16]), .Y(n66) );
endmodule


module CONT ( clk, reset, im_a, im_wen_n, cr_a, curr_time, fb_addr, photo_num, 
        curr_photo_addr, curr_photo_size, en_si, en_init_time, en_fb_addr, 
        en_photo_num, en_curr_photo_addr, en_curr_photo_size, en_so, si_sel, 
        init_time_mux_sel, sftr_n, so_mux_sel, expand_sel );
  output [19:0] im_a;
  output [8:0] cr_a;
  input [23:0] curr_time;
  input [19:0] fb_addr;
  input [1:0] photo_num;
  input [19:0] curr_photo_addr;
  input [1:0] curr_photo_size;
  output [1:0] sftr_n;
  output [1:0] so_mux_sel;
  output [3:0] expand_sel;
  input clk, reset;
  output im_wen_n, en_si, en_init_time, en_fb_addr, en_photo_num,
         en_curr_photo_addr, en_curr_photo_size, en_so, si_sel,
         init_time_mux_sel;
  wire   n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, N138, N139,
         N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, N156, N157, N159, N160, N161, N162,
         N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, N173,
         N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, N184,
         N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, N195,
         N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, N234,
         N235, N236, N237, N238, N239, N240, N241, N242, N243, N266, N267,
         N268, N269, N270, N271, N272, N273, N274, N275, N276, N277, N278,
         N279, N280, N281, N282, N283, N284, N285, N351, N352, N353, N354,
         N355, N356, N357, N358, N359, N390, N391, N392, N393, N394, N395,
         N396, N397, N398, N399, N400, N401, N402, N403, N404, N405, N406,
         N407, N408, N409, N22, N23, N24, N569, N570, N571, N572, N573, N574,
         N575, N576, N577, N590, N591, N592, N593, N594, N595, N608, N609,
         N610, N611, N612, N613, N626, N627, N628, N629, N630, N631, N644,
         N645, N646, N647, N648, N649, N662, N663, N664, N665, N666, N667,
         N671, N676, N719, N720, N721, N722, N723, N724, N725, N726, N727,
         N728, N729, N730, N731, N732, N64, N65, N66, N772, N773, N774, N775,
         N776, N777, N778, N779, N780, N781, N782, N783, N784, N785, N786,
         N787, N788, N789, N790, N791, N795, N796, N797, N798, N799, N800,
         N801, N802, N803, N804, N805, N806, N807, N808, N809, N810, N811,
         N974, N975, N976, N977, N978, N979, N980, N981, N982, N983, N984,
         N985, N986, N987, N988, N989, N990, N991, N992, N993, N994, N995,
         N996, N997, N998, N999, N1000, N1001, N1002, N1003, N1004, N1005,
         N1006, N1007, N1008, N1009, N1010, N1011, N1012, N1013, N1028, N1029,
         N1030, N1031, N1032, N1033, N1034, N1035, N1036, N1037, N1038, N1039,
         N1040, N1041, N1042, N1043, N1044, N1045, N1046, N73, N74, N75, N1062,
         N1063, N1064, N1065, N1066, N1067, N1068, N1069, N1070, N1071, N1072,
         N1073, N1074, N1075, N1076, N1077, N1078, N1079, N1080, N1081, N76,
         N77, N78, N79, N1104, N1105, N1106, N1107, N1108, N1109, N1110, N1111,
         N1112, N1113, N1114, N1115, N1116, N1117, N1118, N1119, N1120, N1121,
         N1122, N80, N81, N82, next_en_si, N1170, N86, N87, N88, N89, N90, N91,
         N1198, N1200, N1201, N1202, N1203, N1204, N1205, N1206, N1207, N1208,
         N1209, N1210, N1211, N1212, N1213, N1214, N1215, N1216, N1217, N1218,
         N1219, N92, N93, N94, N95, _4_net_, _6_net_, N1425, N1447, N1467,
         n378, n379, n420, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         N568, N567, N566, N565, N564, N563, N586, N585, N584, N583, N582,
         N581, N604, N603, N602, N601, N600, N599, N622, N621, N620, N619,
         N618, N617, N640, N639, N638, N637, N636, N635, N658, N657, N656,
         N655, N654, N653, N704, N703, N702, N701, N700, N699, N698, N697,
         N696, N695, N694, N693, N692, \gt_357/A[0] , \add_298/carry[3] ,
         \add_0_root_add_296_2/carry[16] , \add_0_root_add_296_2/carry[15] ,
         \add_0_root_add_296_2/carry[14] , \add_0_root_add_296_2/carry[12] ,
         \add_0_root_add_296_2/carry[8] , \add_0_root_add_296_2/carry[5] ,
         \r864/carry[4] , \r864/carry[5] , \r864/carry[6] , \r864/carry[7] ,
         \r864/carry[8] , \r864/carry[9] , \r864/carry[10] , \r864/carry[11] ,
         \r864/carry[12] , \r864/carry[13] , \r864/carry[14] ,
         \r864/carry[15] , \r864/carry[16] , \r864/carry[17] ,
         \r864/carry[18] , \r864/carry[19] , \sub_358/carry[2] ,
         \sub_358/carry[3] , \sub_358/carry[4] , \sub_358/carry[6] ,
         \sub_358/carry[7] , \sub_358/carry[8] , \sub_358/carry[9] ,
         \sub_358/carry[10] , \sub_358/carry[11] , \sub_358/carry[12] ,
         \sub_358/carry[13] , \sub_358/carry[14] , \sub_358/carry[15] ,
         \sub_358/carry[16] , \sub_358/carry[17] , \sub_358/carry[18] ,
         \sub_358/carry[19] , \r902/carry[19] , \r902/carry[18] ,
         \r902/carry[17] , \r902/carry[16] , \r902/carry[15] ,
         \r902/carry[14] , \r902/carry[13] , \r902/carry[12] ,
         \r902/carry[11] , \r902/carry[10] , \r902/carry[9] , \r902/carry[8] ,
         \r902/carry[7] , \r902/carry[6] , \r902/carry[5] , \r902/carry[4] ,
         \sub_309/carry[4] , \sub_309/carry[5] , \sub_309/carry[6] ,
         \sub_309/carry[7] , \sub_309/carry[8] , \sub_309/carry[9] ,
         \sub_309/carry[10] , \sub_309/carry[11] , \sub_309/carry[12] ,
         \sub_309/carry[13] , \sub_309/carry[14] , \sub_309/carry[15] ,
         \sub_309/carry[16] , \sub_309/carry[17] , \sub_309/carry[18] ,
         \sub_309/carry[19] , \r898/carry[19] , \r898/carry[18] ,
         \r898/carry[17] , \r898/carry[16] , \r898/carry[15] ,
         \r898/carry[14] , \r898/carry[13] , \r898/carry[12] ,
         \r898/carry[11] , \r898/carry[10] , \r898/carry[9] , \r898/carry[8] ,
         \r898/carry[7] , \r898/carry[6] , \add_237/carry[5] , \mult_237/n4 ,
         \mult_237/n3 , \mult_237/n2 , \add_236/carry[5] , \mult_236/n4 ,
         \mult_236/n3 , \mult_236/n2 , \add_235/carry[5] , \mult_235/n4 ,
         \mult_235/n3 , \mult_235/n2 , \add_234/carry[5] , \mult_234/n4 ,
         \mult_234/n3 , \mult_234/n2 , \add_233/carry[5] , \mult_233/n4 ,
         \mult_233/n3 , \mult_233/n2 , \add_232/carry[5] , \mult_232/n4 ,
         \mult_232/n3 , \mult_232/n2 ,
         \add_0_root_add_0_root_add_269_2/carry[2] ,
         \add_0_root_add_0_root_add_269_2/carry[3] ,
         \add_0_root_add_0_root_add_269_2/carry[4] ,
         \add_0_root_add_0_root_add_269_2/carry[9] ,
         \add_0_root_add_0_root_add_269_2/carry[10] ,
         \add_0_root_add_0_root_add_269_2/carry[11] ,
         \add_0_root_add_0_root_add_269_2/carry[12] ,
         \add_0_root_add_0_root_add_269_2/A[0] ,
         \add_0_root_add_0_root_add_269_2/A[1] ,
         \add_0_root_add_0_root_add_269_2/A[2] ,
         \add_0_root_add_0_root_add_269_2/A[3] ,
         \add_0_root_add_0_root_add_269_2/A[8] ,
         \add_0_root_add_0_root_add_269_2/A[9] ,
         \add_0_root_add_0_root_add_269_2/A[10] ,
         \add_0_root_add_0_root_add_269_2/A[11] ,
         \add_0_root_add_0_root_add_269_2/A[12] , \mult_269_2/n26 ,
         \mult_269_2/n25 , \mult_269_2/n24 , \mult_269_2/n23 ,
         \mult_269_2/n22 , \mult_269_2/n21 , \mult_269_2/n20 ,
         \mult_269_2/n19 , \mult_269_2/n18 , \mult_269_2/n17 ,
         \mult_269_2/n16 , \mult_269_2/n15 , \mult_269_2/n14 ,
         \mult_269_2/n13 , \mult_269_2/n12 , \mult_269_2/n11 ,
         \mult_269_2/n10 , \mult_269_2/n9 , \mult_269_2/n8 , \mult_269_2/n7 ,
         \mult_269_2/n6 , \mult_269_2/n5 , \mult_269_2/n4 , \mult_269_2/n3 ,
         \mult_269_2/n2 , n4, n5, n6, n7, n8, n13, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n44, n45, n46, n47, n48,
         n49, n51, n53, n55, n57, n59, n61, n63, n65, n67, n69, n71, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588;
  wire   [2:0] next_state;
  wire   [2:0] state;
  wire   [19:0] work_cntr;
  wire   [19:0] next_work_cntr;
  wire   [19:0] global_cntr;
  wire   [19:0] next_glb_cntr;
  wire   [19:0] write_cntr;
  wire   [8:0] cr_x;
  wire   [19:0] next_write_cntr;
  wire   [8:0] next_cr_x;
  wire   [3:0] h_1;
  wire   [3:0] h_0;
  wire   [3:0] m_1;
  wire   [3:0] m_0;
  wire   [3:0] s_1;
  wire   [3:0] s_0;
  wire   [19:0] read_cntr;
  wire   [8:0] cr_read_cntr;
  wire   [19:0] write_addr;
  wire   [19:0] next_write_addr;
  wire   [1:0] curr_photo;
  wire   [19:0] next_read_cntr;
  wire   [8:0] next_cr_read_cntr;
  wire   [19:0] read_addr;
  wire   [1:0] next_photo;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38;
  assign en_init_time = N1425;
  assign en_curr_photo_addr = N1447;
  assign en_curr_photo_size = N1467;
  assign sftr_n[0] = 1'b0;
  assign sftr_n[1] = 1'b1;

  p_dff_WORD20_NSEL5_0 write_addr_reg ( .clk(clk), .reset(reset), .en(_6_net_), 
        .sel({1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .d(next_write_addr), .q(
        write_addr) );
  p_dff_WORD20_NSEL5_4 read_cntr_reg ( .clk(clk), .reset(reset), .en(_4_net_), 
        .sel({1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .d(next_read_cntr), .q(read_cntr) );
  p_dff_WORD9_NSEL4 cr_read_cntr_reg ( .clk(clk), .reset(reset), .en(_4_net_), 
        .sel({1'b1, 1'b1, 1'b1, 1'b1}), .d(next_cr_read_cntr), .q(cr_read_cntr) );
  p_dff_WORD20_NSEL5_3 write_cntr_reg ( .clk(clk), .reset(reset), .en(_6_net_), 
        .sel({1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .d({n30, n35, n38, 
        next_write_cntr[16:13], n40, next_write_cntr[11:10], n44, 
        next_write_cntr[8:5], n48, next_write_cntr[3:0]}), .q(write_cntr) );
  CONT_DW_div_uns_0 rem_269 ( .a({next_write_cntr[19], n35, n38, 
        next_write_cntr[16:13], n41, next_write_cntr[11:10], n45, 
        next_write_cntr[8:5], n47, next_write_cntr[3], n32, next_write_cntr[1], 
        n27}), .b({1'b1, 1'b1, 1'b0, 1'b1}), .remainder({
        \add_0_root_add_0_root_add_269_2/A[3] , 
        \add_0_root_add_0_root_add_269_2/A[2] , 
        \add_0_root_add_0_root_add_269_2/A[1] , 
        \add_0_root_add_0_root_add_269_2/A[0] }) );
  CONT_DW01_inc_0 add_192 ( .A({1'b0, cr_read_cntr}), .SUM({
        SYNOPSYS_UNCONNECTED__0, N359, N358, N357, N356, N355, N354, N353, 
        N352, N351}) );
  CONT_DW01_inc_1 add_185 ( .A({1'b0, read_cntr}), .SUM({
        SYNOPSYS_UNCONNECTED__1, N243, N242, N241, N240, N239, N238, N237, 
        N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, 
        N224}) );
  CONT_DW_div_uns_1 rem_153 ( .a(curr_time[7:0]), .b({1'b1, 1'b0, 1'b1, 1'b0}), 
        .remainder({s_0[3:1], N653}) );
  CONT_DW_div_uns_2 div_152 ( .a(curr_time[7:0]), .b({1'b1, 1'b0, 1'b1, 1'b0}), 
        .quotient({SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, s_1[3:1], N635}) );
  CONT_DW_div_uns_3 rem_151 ( .a(curr_time[15:8]), .b({1'b1, 1'b0, 1'b1, 1'b0}), .remainder({m_0[3:1], N617}) );
  CONT_DW_div_uns_4 div_150 ( .a(curr_time[15:8]), .b({1'b1, 1'b0, 1'b1, 1'b0}), .quotient({SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, m_1[3:1], N599}) );
  CONT_DW_div_uns_5 rem_149 ( .a(curr_time[23:16]), .b({1'b1, 1'b0, 1'b1, 1'b0}), .remainder({h_0[3:1], N581}) );
  CONT_DW_div_uns_6 div_148 ( .a(curr_time[23:16]), .b({1'b1, 1'b0, 1'b1, 1'b0}), .quotient({SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, h_1[3:1], N563})
         );
  CONT_DW_div_uns_8 div_146 ( .a({n30, next_write_cntr[18:3], n33, 
        next_write_cntr[1:0]}), .b({1'b1, 1'b1, 1'b0, 1'b1}), .quotient({
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, N195, N194, N193, N192, N191, N190, N189, 
        N188, N187, N186, N185, N184, N183, N182, N181, N180, N179}) );
  CONT_DW_div_uns_9 div_145 ( .a({n29, n35, n37, next_write_cntr[16:13], n40, 
        next_write_cntr[11:10], n44, next_write_cntr[8:5], n48, 
        next_write_cntr[3], n33, next_write_cntr[1:0]}), .b({1'b1, 1'b0, 1'b0, 
        1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0}), .quotient({
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24, 
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, next_cr_x[8:2], N693, N692}) );
  CONT_DW01_add_33 r889 ( .A(write_addr), .B(fb_addr), .CI(1'b0), .SUM({N811, 
        N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, 
        N798, N797, N796, N795, N976, N975, N974}) );
  CONT_DW01_add_34 r888 ( .A(read_addr), .B(curr_photo_addr), .CI(1'b0), .SUM(
        {N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, 
        N780, N779, N778, N777, N776, N775, N774, N773, N772}) );
  CONT_DW_div_uns_11 div_142 ( .a(write_cntr), .b({1'b1, 1'b0, 1'b0, 1'b1, 
        1'b1, 1'b1, 1'b0, 1'b0, 1'b0}), .quotient({SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, 
        SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, SYNOPSYS_UNCONNECTED__34, 
        SYNOPSYS_UNCONNECTED__35, SYNOPSYS_UNCONNECTED__36, 
        SYNOPSYS_UNCONNECTED__37, SYNOPSYS_UNCONNECTED__38, cr_x}) );
  CONT_DW_div_uns_12 r865 ( .a({n8, n8, n8, n8, n8, n8, n8, n8, n8, n8, n8, n8, 
        N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, 
        N397, N396, N395, N394, N393, N392, N391, N390}), .b({1'b1, 1'b1, 1'b0}), .remainder({N24, N23, N22}) );
  CONT_DW_div_uns_13 rem_358 ( .a({n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, 
        n7, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, 
        N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, 
        N1200}), .b({1'b1, 1'b1, 1'b1, 1'b0}), .remainder({N95, N94, N93, N92}) );
  CONT_DW_div_uns_14 rem_353_2 ( .a({N1170, N157, N156, N155, N154, N153, N152, 
        N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, 
        N139, N138}), .b({1'b1, 1'b0, 1'b1}), .remainder({N91, N90, N89}) );
  CONT_DW_div_uns_15 rem_353 ( .a({N1170, N157, N156, N155, N154, N153, N152, 
        N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, 
        N139, N138}), .b({1'b1, 1'b0, 1'b1}), .remainder({N88, N87, N86}) );
  CONT_DW_div_uns_16 r903 ( .a({n6, n6, n6, n6, n6, n6, n6, n6, n6, n6, n6, n6, 
        N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, 
        N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, n219}), 
        .b({1'b1, 1'b1, 1'b0}), .remainder({N82, N81, N80}) );
  CONT_DW01_inc_2 r860 ( .A(write_cntr), .SUM({N285, N284, N283, N282, N281, 
        N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, 
        N268, N267, N266}) );
  CONT_DW01_inc_3 r842 ( .A({1'b0, n85, n74, work_cntr[17], n79, n94, n90, n81, 
        n92, n87, n77, n102, n98, n100, n96, n83, work_cntr[4], n218, n217, 
        n216, n219}), .SUM({N1170, N157, N156, N155, N154, N153, N152, N151, 
        N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, 
        N138}) );
  CONT_DW_div_uns_17 r885 ( .a({n85, n74, work_cntr[17], n79, n94, n90, n81, 
        n92, n88, n76, n102, n98, n100, n96, n83, work_cntr[4], n218, n217, 
        n216, n219}), .b({1'b1, 1'b0, 1'b1}), .remainder({N66, N65, N64}) );
  CONT_DW_div_uns_18 rem_309 ( .a({n5, n5, n5, n5, n5, n5, n5, n5, n5, n5, n5, 
        n5, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, 
        N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, 
        N390}), .b({1'b1, 1'b1, 1'b0}), .remainder({N75, N74, N73}) );
  CONT_DW01_inc_4 add_130 ( .A({global_cntr[19:1], N994}), .SUM({N178, N177, 
        N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, 
        N164, N163, N162, N161, N160, N159}) );
  CONT_DW_div_uns_19 r899 ( .a({n4, n4, n4, n4, n4, n4, n4, n4, n4, n4, n4, n4, 
        N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, 
        N1071, N1070, N1069, N1068, N1067, N1066, n218, n217, n216, n219}), 
        .b({1'b1, 1'b1, 1'b1, 1'b0}), .remainder({N79, N78, N77, N76}) );
  ADDHXL \mult_237/U5  ( .A(N653), .B(s_0[1]), .CO(\mult_237/n4 ), .S(N654) );
  ADDFXL \mult_237/U4  ( .A(s_0[2]), .B(s_0[1]), .CI(\mult_237/n4 ), .CO(
        \mult_237/n3 ), .S(N655) );
  ADDFXL \mult_237/U3  ( .A(s_0[3]), .B(s_0[2]), .CI(\mult_237/n3 ), .CO(
        \mult_237/n2 ), .S(N656) );
  ADDHXL \mult_236/U5  ( .A(N635), .B(s_1[1]), .CO(\mult_236/n4 ), .S(N636) );
  ADDFXL \mult_236/U4  ( .A(s_1[2]), .B(s_1[1]), .CI(\mult_236/n4 ), .CO(
        \mult_236/n3 ), .S(N637) );
  ADDFXL \mult_236/U3  ( .A(s_1[3]), .B(s_1[2]), .CI(\mult_236/n3 ), .CO(
        \mult_236/n2 ), .S(N638) );
  ADDHXL \mult_235/U5  ( .A(N617), .B(m_0[1]), .CO(\mult_235/n4 ), .S(N618) );
  ADDFXL \mult_235/U4  ( .A(m_0[2]), .B(m_0[1]), .CI(\mult_235/n4 ), .CO(
        \mult_235/n3 ), .S(N619) );
  ADDFXL \mult_235/U3  ( .A(m_0[3]), .B(m_0[2]), .CI(\mult_235/n3 ), .CO(
        \mult_235/n2 ), .S(N620) );
  ADDHXL \mult_234/U5  ( .A(N599), .B(m_1[1]), .CO(\mult_234/n4 ), .S(N600) );
  ADDFXL \mult_234/U4  ( .A(m_1[2]), .B(m_1[1]), .CI(\mult_234/n4 ), .CO(
        \mult_234/n3 ), .S(N601) );
  ADDFXL \mult_234/U3  ( .A(m_1[3]), .B(m_1[2]), .CI(\mult_234/n3 ), .CO(
        \mult_234/n2 ), .S(N602) );
  ADDHXL \mult_233/U5  ( .A(N581), .B(h_0[1]), .CO(\mult_233/n4 ), .S(N582) );
  ADDFXL \mult_233/U4  ( .A(h_0[2]), .B(h_0[1]), .CI(\mult_233/n4 ), .CO(
        \mult_233/n3 ), .S(N583) );
  ADDFXL \mult_233/U3  ( .A(h_0[3]), .B(h_0[2]), .CI(\mult_233/n3 ), .CO(
        \mult_233/n2 ), .S(N584) );
  ADDHXL \mult_232/U5  ( .A(N563), .B(h_1[1]), .CO(\mult_232/n4 ), .S(N564) );
  ADDFXL \mult_232/U4  ( .A(h_1[2]), .B(h_1[1]), .CI(\mult_232/n4 ), .CO(
        \mult_232/n3 ), .S(N565) );
  ADDFXL \mult_232/U3  ( .A(h_1[3]), .B(h_1[2]), .CI(\mult_232/n3 ), .CO(
        \mult_232/n2 ), .S(N566) );
  ADDHXL \mult_269_2/U19  ( .A(next_cr_x[3]), .B(N693), .CO(\mult_269_2/n25 ), 
        .S(\mult_269_2/n26 ) );
  ADDFXL \mult_269_2/U18  ( .A(N693), .B(next_cr_x[4]), .CI(next_cr_x[2]), 
        .CO(\mult_269_2/n23 ), .S(\mult_269_2/n24 ) );
  ADDFXL \mult_269_2/U17  ( .A(next_cr_x[2]), .B(next_cr_x[5]), .CI(
        next_cr_x[3]), .CO(\mult_269_2/n21 ), .S(\mult_269_2/n22 ) );
  ADDFXL \mult_269_2/U16  ( .A(next_cr_x[3]), .B(next_cr_x[6]), .CI(
        next_cr_x[4]), .CO(\mult_269_2/n19 ), .S(\mult_269_2/n20 ) );
  ADDFXL \mult_269_2/U15  ( .A(next_cr_x[4]), .B(next_cr_x[7]), .CI(
        next_cr_x[5]), .CO(\mult_269_2/n17 ), .S(\mult_269_2/n18 ) );
  ADDFXL \mult_269_2/U14  ( .A(next_cr_x[5]), .B(next_cr_x[8]), .CI(
        next_cr_x[6]), .CO(\mult_269_2/n15 ), .S(\mult_269_2/n16 ) );
  ADDHXL \mult_269_2/U13  ( .A(next_cr_x[7]), .B(next_cr_x[6]), .CO(
        \mult_269_2/n13 ), .S(\mult_269_2/n14 ) );
  ADDHXL \mult_269_2/U12  ( .A(next_cr_x[8]), .B(next_cr_x[7]), .CO(
        \mult_269_2/n11 ), .S(\mult_269_2/n12 ) );
  ADDHXL \mult_269_2/U11  ( .A(N692), .B(next_cr_x[2]), .CO(\mult_269_2/n10 ), 
        .S(N694) );
  ADDFXL \mult_269_2/U10  ( .A(\mult_269_2/n10 ), .B(N692), .CI(
        \mult_269_2/n26 ), .CO(\mult_269_2/n9 ), .S(N695) );
  ADDFXL \mult_269_2/U9  ( .A(\mult_269_2/n24 ), .B(\mult_269_2/n25 ), .CI(
        \mult_269_2/n9 ), .CO(\mult_269_2/n8 ), .S(N696) );
  ADDFXL \mult_269_2/U8  ( .A(\mult_269_2/n22 ), .B(\mult_269_2/n23 ), .CI(
        \mult_269_2/n8 ), .CO(\mult_269_2/n7 ), .S(N697) );
  ADDFXL \mult_269_2/U7  ( .A(\mult_269_2/n20 ), .B(\mult_269_2/n21 ), .CI(
        \mult_269_2/n7 ), .CO(\mult_269_2/n6 ), .S(N698) );
  ADDFXL \mult_269_2/U6  ( .A(\mult_269_2/n18 ), .B(\mult_269_2/n19 ), .CI(
        \mult_269_2/n6 ), .CO(\mult_269_2/n5 ), .S(N699) );
  ADDFXL \mult_269_2/U5  ( .A(\mult_269_2/n16 ), .B(\mult_269_2/n17 ), .CI(
        \mult_269_2/n5 ), .CO(\mult_269_2/n4 ), .S(N700) );
  ADDFXL \mult_269_2/U4  ( .A(\mult_269_2/n15 ), .B(\mult_269_2/n14 ), .CI(
        \mult_269_2/n4 ), .CO(\mult_269_2/n3 ), .S(N701) );
  ADDFXL \mult_269_2/U3  ( .A(\mult_269_2/n12 ), .B(\mult_269_2/n13 ), .CI(
        \mult_269_2/n3 ), .CO(\mult_269_2/n2 ), .S(N702) );
  ADDFXL \mult_269_2/U2  ( .A(\mult_269_2/n11 ), .B(next_cr_x[8]), .CI(
        \mult_269_2/n2 ), .CO(N704), .S(N703) );
  CONT_DW_div_uns_59 r868 ( .a(cr_read_cntr), .b({1'b1, 1'b1, 1'b0, 1'b0, 1'b0}), .remainder({N676, N671, N571, N570, N569}) );
  CONT_DW_div_uns_71 rem_146 ( .a({1'b0, 1'b0, 1'b0, N195, N194, N193, N192, 
        N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, 
        N179}), .b({1'b1, 1'b1, 1'b0, 1'b0, 1'b0}), .remainder({
        \add_0_root_add_0_root_add_269_2/A[12] , 
        \add_0_root_add_0_root_add_269_2/A[11] , 
        \add_0_root_add_0_root_add_269_2/A[10] , 
        \add_0_root_add_0_root_add_269_2/A[9] , 
        \add_0_root_add_0_root_add_269_2/A[8] }) );
  DFFSX1 en_si_reg ( .D(next_en_si), .CK(clk), .SN(n588), .Q(en_si) );
  ADDFXL \add_298/U1_2  ( .A(global_cntr[2]), .B(curr_photo[1]), .CI(n25), 
        .CO(\add_298/carry[3] ), .S(N996) );
  ADDFXL \add_0_root_add_0_root_add_269_2/U1_1  ( .A(
        \add_0_root_add_0_root_add_269_2/A[1] ), .B(N693), .CI(n16), .CO(
        \add_0_root_add_0_root_add_269_2/carry[2] ), .S(N720) );
  ADDFXL \add_0_root_add_0_root_add_269_2/U1_2  ( .A(
        \add_0_root_add_0_root_add_269_2/A[2] ), .B(N694), .CI(
        \add_0_root_add_0_root_add_269_2/carry[2] ), .CO(
        \add_0_root_add_0_root_add_269_2/carry[3] ), .S(N721) );
  ADDFXL \add_0_root_add_0_root_add_269_2/U1_3  ( .A(
        \add_0_root_add_0_root_add_269_2/A[3] ), .B(N695), .CI(
        \add_0_root_add_0_root_add_269_2/carry[3] ), .CO(
        \add_0_root_add_0_root_add_269_2/carry[4] ), .S(N722) );
  ADDFXL \add_0_root_add_0_root_add_269_2/U1_8  ( .A(
        \add_0_root_add_0_root_add_269_2/A[8] ), .B(N700), .CI(n15), .CO(
        \add_0_root_add_0_root_add_269_2/carry[9] ), .S(N727) );
  ADDFXL \add_0_root_add_0_root_add_269_2/U1_9  ( .A(
        \add_0_root_add_0_root_add_269_2/A[9] ), .B(N701), .CI(
        \add_0_root_add_0_root_add_269_2/carry[9] ), .CO(
        \add_0_root_add_0_root_add_269_2/carry[10] ), .S(N728) );
  ADDFXL \add_0_root_add_0_root_add_269_2/U1_12  ( .A(
        \add_0_root_add_0_root_add_269_2/A[12] ), .B(N704), .CI(
        \add_0_root_add_0_root_add_269_2/carry[12] ), .CO(N732), .S(N731) );
  ADDFXL \add_0_root_add_0_root_add_269_2/U1_11  ( .A(
        \add_0_root_add_0_root_add_269_2/A[11] ), .B(N703), .CI(
        \add_0_root_add_0_root_add_269_2/carry[11] ), .CO(
        \add_0_root_add_0_root_add_269_2/carry[12] ), .S(N730) );
  ADDFXL \add_0_root_add_0_root_add_269_2/U1_10  ( .A(
        \add_0_root_add_0_root_add_269_2/A[10] ), .B(N702), .CI(
        \add_0_root_add_0_root_add_269_2/carry[10] ), .CO(
        \add_0_root_add_0_root_add_269_2/carry[11] ), .S(N729) );
  ADDFXL \add_237/U1_4  ( .A(N654), .B(N676), .CI(n24), .CO(\add_237/carry[5] ), .S(N663) );
  ADDFXL \add_235/U1_4  ( .A(N618), .B(N676), .CI(n23), .CO(\add_235/carry[5] ), .S(N627) );
  ADDFXL \add_233/U1_4  ( .A(N582), .B(N676), .CI(n22), .CO(\add_233/carry[5] ), .S(N591) );
  ADDFXL \add_236/U1_4  ( .A(N636), .B(N676), .CI(n21), .CO(\add_236/carry[5] ), .S(N645) );
  ADDFXL \add_234/U1_4  ( .A(N600), .B(N676), .CI(n20), .CO(\add_234/carry[5] ), .S(N609) );
  ADDFXL \add_232/U1_4  ( .A(N564), .B(N676), .CI(n19), .CO(\add_232/carry[5] ), .S(N573) );
  DFFRHQX1 \state_reg[2]  ( .D(n573), .CK(clk), .RN(n588), .Q(state[2]) );
  DFFRHQX1 \state_reg[0]  ( .D(next_state[0]), .CK(clk), .RN(n588), .Q(
        state[0]) );
  DFFRHQX1 \work_cntr_reg[13]  ( .D(next_work_cntr[13]), .CK(clk), .RN(n588), 
        .Q(work_cntr[13]) );
  DFFRHQX1 \work_cntr_reg[15]  ( .D(next_work_cntr[15]), .CK(clk), .RN(n588), 
        .Q(work_cntr[15]) );
  DFFRHQX1 \work_cntr_reg[14]  ( .D(next_work_cntr[14]), .CK(clk), .RN(n588), 
        .Q(work_cntr[14]) );
  DFFRHQX1 \work_cntr_reg[11]  ( .D(next_work_cntr[11]), .CK(clk), .RN(n588), 
        .Q(work_cntr[11]) );
  DFFRHQX1 \work_cntr_reg[16]  ( .D(next_work_cntr[16]), .CK(clk), .RN(n588), 
        .Q(work_cntr[16]) );
  DFFRHQX1 \work_cntr_reg[12]  ( .D(next_work_cntr[12]), .CK(clk), .RN(n588), 
        .Q(work_cntr[12]) );
  DFFRHQX1 \work_cntr_reg[8]  ( .D(next_work_cntr[8]), .CK(clk), .RN(n588), 
        .Q(work_cntr[8]) );
  DFFRHQX1 \work_cntr_reg[9]  ( .D(next_work_cntr[9]), .CK(clk), .RN(n588), 
        .Q(work_cntr[9]) );
  DFFRHQX1 \work_cntr_reg[10]  ( .D(next_work_cntr[10]), .CK(clk), .RN(n588), 
        .Q(work_cntr[10]) );
  DFFRHQX1 \work_cntr_reg[5]  ( .D(next_work_cntr[5]), .CK(clk), .RN(n588), 
        .Q(work_cntr[5]) );
  DFFRHQX1 \work_cntr_reg[6]  ( .D(next_work_cntr[6]), .CK(clk), .RN(n588), 
        .Q(work_cntr[6]) );
  DFFRHQX1 \work_cntr_reg[7]  ( .D(next_work_cntr[7]), .CK(clk), .RN(n588), 
        .Q(work_cntr[7]) );
  DFFRHQX1 \work_cntr_reg[18]  ( .D(next_work_cntr[18]), .CK(clk), .RN(n588), 
        .Q(work_cntr[18]) );
  DFFRHQX1 \work_cntr_reg[19]  ( .D(next_work_cntr[19]), .CK(clk), .RN(n588), 
        .Q(work_cntr[19]) );
  DFFRHQX1 \work_cntr_reg[3]  ( .D(next_work_cntr[3]), .CK(clk), .RN(n588), 
        .Q(N1065) );
  DFFRHQX1 \work_cntr_reg[0]  ( .D(\gt_357/A[0] ), .CK(clk), .RN(n588), .Q(
        N1062) );
  DFFRHQX1 \work_cntr_reg[2]  ( .D(next_work_cntr[2]), .CK(clk), .RN(n588), 
        .Q(N1064) );
  DFFRHQX1 \work_cntr_reg[1]  ( .D(next_work_cntr[1]), .CK(clk), .RN(n588), 
        .Q(N1063) );
  DFFSRX1 \global_cntr_reg[3]  ( .D(n586), .CK(clk), .SN(1'b1), .RN(n588), .Q(
        global_cntr[3]), .QN(n452) );
  DFFSRX1 \global_cntr_reg[4]  ( .D(n585), .CK(clk), .SN(1'b1), .RN(n588), .Q(
        global_cntr[4]), .QN(n451) );
  DFFSRX1 \global_cntr_reg[0]  ( .D(next_glb_cntr[0]), .CK(clk), .SN(1'b1), 
        .RN(n588), .Q(N994), .QN(n455) );
  DFFSRX1 \global_cntr_reg[5]  ( .D(next_glb_cntr[5]), .CK(clk), .SN(1'b1), 
        .RN(n588), .Q(global_cntr[5]), .QN(n450) );
  DFFSRX1 \global_cntr_reg[6]  ( .D(next_glb_cntr[6]), .CK(clk), .SN(1'b1), 
        .RN(n588), .Q(global_cntr[6]), .QN(n449) );
  DFFSRX1 \global_cntr_reg[7]  ( .D(n584), .CK(clk), .SN(1'b1), .RN(n588), .Q(
        global_cntr[7]), .QN(n448) );
  DFFSRX1 \global_cntr_reg[8]  ( .D(n583), .CK(clk), .SN(1'b1), .RN(n588), .Q(
        global_cntr[8]), .QN(n447) );
  DFFSRX1 \global_cntr_reg[9]  ( .D(n582), .CK(clk), .SN(1'b1), .RN(n588), .Q(
        global_cntr[9]), .QN(n446) );
  DFFSRX1 \global_cntr_reg[10]  ( .D(n581), .CK(clk), .SN(1'b1), .RN(n588), 
        .Q(global_cntr[10]), .QN(n445) );
  DFFSRX1 \global_cntr_reg[11]  ( .D(n580), .CK(clk), .SN(1'b1), .RN(n588), 
        .Q(global_cntr[11]), .QN(n444) );
  DFFSRX1 \global_cntr_reg[12]  ( .D(n579), .CK(clk), .SN(1'b1), .RN(n588), 
        .Q(global_cntr[12]), .QN(n443) );
  DFFSRX1 \global_cntr_reg[13]  ( .D(n578), .CK(clk), .SN(1'b1), .RN(n588), 
        .Q(global_cntr[13]), .QN(n442) );
  DFFSRX1 \global_cntr_reg[14]  ( .D(next_glb_cntr[14]), .CK(clk), .SN(1'b1), 
        .RN(n588), .Q(global_cntr[14]), .QN(n441) );
  DFFSRX1 \global_cntr_reg[15]  ( .D(next_glb_cntr[15]), .CK(clk), .SN(1'b1), 
        .RN(n588), .Q(global_cntr[15]), .QN(n440) );
  DFFSRX1 \global_cntr_reg[16]  ( .D(n577), .CK(clk), .SN(1'b1), .RN(n588), 
        .Q(global_cntr[16]), .QN(n439) );
  DFFSRX1 \global_cntr_reg[17]  ( .D(n576), .CK(clk), .SN(1'b1), .RN(n588), 
        .Q(global_cntr[17]), .QN(n438) );
  DFFSRX1 \global_cntr_reg[18]  ( .D(n575), .CK(clk), .SN(1'b1), .RN(n588), 
        .Q(global_cntr[18]), .QN(n437) );
  DFFSRX1 \global_cntr_reg[19]  ( .D(n574), .CK(clk), .SN(1'b1), .RN(n588), 
        .Q(global_cntr[19]), .QN(n420) );
  DFFSRX1 \curr_photo_reg[0]  ( .D(next_photo[0]), .CK(clk), .SN(1'b1), .RN(
        n588), .Q(curr_photo[0]), .QN(n379) );
  DFFSRX1 \curr_photo_reg[1]  ( .D(next_photo[1]), .CK(clk), .SN(1'b1), .RN(
        n588), .Q(curr_photo[1]), .QN(n378) );
  DFFRHQX4 \work_cntr_reg[17]  ( .D(next_work_cntr[17]), .CK(clk), .RN(n588), 
        .Q(work_cntr[17]) );
  DFFRX2 \state_reg[1]  ( .D(next_state[1]), .CK(clk), .RN(n588), .QN(n525) );
  DFFRX2 \global_cntr_reg[2]  ( .D(n587), .CK(clk), .RN(n588), .Q(
        global_cntr[2]), .QN(n453) );
  DFFRX2 \global_cntr_reg[1]  ( .D(next_glb_cntr[1]), .CK(clk), .RN(n588), .Q(
        global_cntr[1]), .QN(n454) );
  DFFRHQX4 \work_cntr_reg[4]  ( .D(next_work_cntr[4]), .CK(clk), .RN(n588), 
        .Q(work_cntr[4]) );
  OAI21X2 U5 ( .A0(state[2]), .A1(n525), .B0(n526), .Y(en_so) );
  AOI221X1 U6 ( .A0(n543), .A1(n214), .B0(n544), .B1(n545), .C0(n503), .Y(n542) );
  NOR2X1 U7 ( .A(n85), .B(\r898/carry[19] ), .Y(n4) );
  NOR2X1 U8 ( .A(work_cntr[19]), .B(\sub_309/carry[19] ), .Y(n5) );
  NOR2XL U9 ( .A(n85), .B(\r902/carry[19] ), .Y(n6) );
  NOR2X1 U10 ( .A(next_work_cntr[19]), .B(\sub_358/carry[19] ), .Y(n7) );
  NOR2X1 U11 ( .A(work_cntr[19]), .B(\r864/carry[19] ), .Y(n8) );
  AND3X2 U12 ( .A(n351), .B(n349), .C(n541), .Y(n13) );
  INVXL U13 ( .A(next_write_cntr[9]), .Y(n42) );
  INVXL U14 ( .A(next_write_cntr[4]), .Y(n46) );
  CLKINVX1 U15 ( .A(n31), .Y(n33) );
  AO22XL U16 ( .A0(write_cntr[2]), .A1(n201), .B0(N268), .B1(n200), .Y(
        next_write_cntr[2]) );
  NAND3X1 U17 ( .A(n525), .B(n536), .C(n414), .Y(init_time_mux_sel) );
  AND2X2 U18 ( .A(N699), .B(n143), .Y(n15) );
  AND2X2 U19 ( .A(N692), .B(\add_0_root_add_0_root_add_269_2/A[0] ), .Y(n16)
         );
  OR2X1 U20 ( .A(n526), .B(state[0]), .Y(n17) );
  OA22X1 U21 ( .A0(n221), .A1(n339), .B0(n328), .B1(n329), .Y(n18) );
  AND2X2 U22 ( .A(N671), .B(N563), .Y(n19) );
  AND2X2 U23 ( .A(N671), .B(N599), .Y(n20) );
  AND2X2 U24 ( .A(N671), .B(N635), .Y(n21) );
  AND2X2 U25 ( .A(N671), .B(N581), .Y(n22) );
  AND2X2 U26 ( .A(N671), .B(N617), .Y(n23) );
  AND2X2 U27 ( .A(N671), .B(N653), .Y(n24) );
  AND2X2 U28 ( .A(curr_photo[0]), .B(global_cntr[1]), .Y(n25) );
  NOR3X2 U29 ( .A(n432), .B(n454), .C(n453), .Y(N1467) );
  NOR2X2 U30 ( .A(n220), .B(n335), .Y(next_work_cntr[2]) );
  NOR2X2 U31 ( .A(n220), .B(n336), .Y(next_work_cntr[1]) );
  NOR2X2 U32 ( .A(n220), .B(n334), .Y(next_work_cntr[4]) );
  INVX3 U33 ( .A(n73), .Y(n74) );
  NOR2BX2 U34 ( .AN(n460), .B(N676), .Y(n467) );
  AND4X2 U35 ( .A(n490), .B(n491), .C(n489), .D(n492), .Y(n460) );
  OAI33X1 U36 ( .A0(n411), .A1(n310), .A2(n309), .B0(n232), .B1(n240), .B2(
        n407), .Y(n410) );
  OAI21X1 U37 ( .A0(N23), .A1(N22), .B0(N24), .Y(n407) );
  ADDHX1 U38 ( .A(h_0[3]), .B(\mult_233/n2 ), .CO(N586), .S(N585) );
  ADDHX1 U39 ( .A(m_0[3]), .B(\mult_235/n2 ), .CO(N622), .S(N621) );
  ADDHX1 U40 ( .A(s_0[3]), .B(\mult_237/n2 ), .CO(N658), .S(N657) );
  NOR4XL U41 ( .A(n455), .B(n454), .C(n453), .D(n452), .Y(n562) );
  AND3XL U42 ( .A(write_cntr[8]), .B(write_cntr[6]), .C(write_cntr[7]), .Y(
        n566) );
  NOR4X4 U43 ( .A(write_cntr[16]), .B(write_cntr[17]), .C(write_cntr[18]), .D(
        write_cntr[19]), .Y(n328) );
  AOI222X4 U48 ( .A0(n213), .A1(next_write_cntr[3]), .B0(write_addr[3]), .B1(
        n199), .C0(N722), .C1(n205), .Y(n266) );
  AOI222X4 U49 ( .A0(n213), .A1(n47), .B0(write_addr[4]), .B1(n199), .C0(N723), 
        .C1(n205), .Y(n263) );
  NOR2X2 U50 ( .A(n412), .B(n309), .Y(n300) );
  AOI32XL U51 ( .A0(n407), .A1(n241), .A2(n300), .B0(n238), .B1(n408), .Y(n406) );
  AOI2BB1X2 U52 ( .A0N(n306), .A1N(n426), .B0(n506), .Y(n238) );
  INVXL U53 ( .A(next_write_cntr[0]), .Y(n26) );
  CLKINVX1 U54 ( .A(n26), .Y(n27) );
  OAI221X1 U55 ( .A0(n230), .A1(n231), .B0(n232), .B1(n233), .C0(n212), .Y(
        so_mux_sel[1]) );
  AOI222X4 U56 ( .A0(n213), .A1(next_write_cntr[5]), .B0(write_addr[5]), .B1(
        n199), .C0(N724), .C1(n205), .Y(n257) );
  MXI2XL U57 ( .A(n505), .B(n238), .S0(n240), .Y(n504) );
  NAND2X1 U58 ( .A(n300), .B(n240), .Y(n231) );
  AOI2BB1X2 U59 ( .A0N(n230), .A1N(n426), .B0(n506), .Y(n240) );
  NOR3XL U60 ( .A(write_cntr[13]), .B(write_cntr[15]), .C(write_cntr[14]), .Y(
        n565) );
  INVXL U61 ( .A(next_write_cntr[19]), .Y(n28) );
  INVXL U62 ( .A(n28), .Y(n29) );
  INVX1 U63 ( .A(n28), .Y(n30) );
  CLKINVX1 U64 ( .A(next_write_cntr[2]), .Y(n31) );
  CLKINVX1 U65 ( .A(n31), .Y(n32) );
  INVX1 U66 ( .A(next_write_cntr[18]), .Y(n34) );
  CLKINVX1 U67 ( .A(n34), .Y(n35) );
  CLKINVX1 U68 ( .A(next_write_cntr[17]), .Y(n36) );
  CLKINVX1 U69 ( .A(n36), .Y(n37) );
  INVX1 U70 ( .A(n36), .Y(n38) );
  CLKINVX1 U71 ( .A(next_write_cntr[12]), .Y(n39) );
  INVXL U72 ( .A(n39), .Y(n40) );
  INVX1 U74 ( .A(n39), .Y(n41) );
  INVXL U75 ( .A(n42), .Y(n44) );
  INVX1 U76 ( .A(n42), .Y(n45) );
  CLKINVX1 U77 ( .A(n46), .Y(n47) );
  INVXL U78 ( .A(n46), .Y(n48) );
  CLKINVX1 U79 ( .A(n591), .Y(n49) );
  INVX16 U80 ( .A(n49), .Y(im_a[19]) );
  CLKINVX1 U81 ( .A(n592), .Y(n51) );
  INVX16 U82 ( .A(n51), .Y(im_a[18]) );
  CLKINVX1 U83 ( .A(n593), .Y(n53) );
  INVX16 U84 ( .A(n53), .Y(im_a[17]) );
  CLKINVX1 U85 ( .A(n594), .Y(n55) );
  INVX16 U86 ( .A(n55), .Y(im_a[16]) );
  CLKINVX1 U87 ( .A(n595), .Y(n57) );
  INVX16 U88 ( .A(n57), .Y(im_a[15]) );
  CLKINVX1 U89 ( .A(n596), .Y(n59) );
  INVX16 U90 ( .A(n59), .Y(im_a[14]) );
  CLKINVX1 U91 ( .A(n597), .Y(n61) );
  INVX16 U92 ( .A(n61), .Y(im_a[13]) );
  CLKINVX1 U93 ( .A(n598), .Y(n63) );
  INVX16 U94 ( .A(n63), .Y(im_a[12]) );
  CLKINVX1 U95 ( .A(n599), .Y(n65) );
  INVX16 U96 ( .A(n65), .Y(im_a[11]) );
  CLKINVX1 U97 ( .A(n600), .Y(n67) );
  INVX16 U98 ( .A(n67), .Y(im_a[10]) );
  INVX1 U99 ( .A(n610), .Y(n69) );
  INVX16 U100 ( .A(n69), .Y(im_a[0]) );
  OAI211XL U101 ( .A0(n455), .A1(n208), .B0(n403), .C0(n404), .Y(n610) );
  CLKINVX1 U102 ( .A(n613), .Y(n71) );
  INVX16 U103 ( .A(n71), .Y(cr_a[7]) );
  CLKINVX1 U104 ( .A(work_cntr[18]), .Y(n73) );
  CLKINVX1 U105 ( .A(work_cntr[10]), .Y(n75) );
  CLKINVX1 U106 ( .A(n75), .Y(n76) );
  CLKINVX1 U107 ( .A(n75), .Y(n77) );
  CLKINVX1 U108 ( .A(work_cntr[16]), .Y(n78) );
  CLKINVX2 U109 ( .A(n78), .Y(n79) );
  CLKINVX1 U110 ( .A(work_cntr[13]), .Y(n80) );
  CLKINVX2 U111 ( .A(n80), .Y(n81) );
  CLKINVX1 U112 ( .A(work_cntr[5]), .Y(n82) );
  INVX3 U113 ( .A(n82), .Y(n83) );
  CLKINVX1 U114 ( .A(work_cntr[19]), .Y(n84) );
  CLKINVX2 U115 ( .A(n84), .Y(n85) );
  CLKINVX1 U116 ( .A(work_cntr[11]), .Y(n86) );
  CLKINVX1 U117 ( .A(n86), .Y(n87) );
  CLKINVX1 U118 ( .A(n86), .Y(n88) );
  CLKINVX1 U119 ( .A(work_cntr[14]), .Y(n89) );
  CLKINVX2 U120 ( .A(n89), .Y(n90) );
  CLKINVX1 U121 ( .A(work_cntr[12]), .Y(n91) );
  CLKINVX2 U122 ( .A(n91), .Y(n92) );
  CLKINVX1 U123 ( .A(work_cntr[15]), .Y(n93) );
  CLKINVX2 U124 ( .A(n93), .Y(n94) );
  CLKINVX1 U125 ( .A(work_cntr[6]), .Y(n95) );
  INVX3 U126 ( .A(n95), .Y(n96) );
  CLKINVX1 U127 ( .A(work_cntr[8]), .Y(n97) );
  INVX3 U128 ( .A(n97), .Y(n98) );
  CLKINVX1 U129 ( .A(work_cntr[7]), .Y(n99) );
  INVX3 U130 ( .A(n99), .Y(n100) );
  CLKINVX1 U131 ( .A(work_cntr[9]), .Y(n101) );
  INVX3 U132 ( .A(n101), .Y(n102) );
  OR2XL U133 ( .A(n83), .B(work_cntr[4]), .Y(\r898/carry[6] ) );
  INVX8 U134 ( .A(reset), .Y(n588) );
  NOR4XL U155 ( .A(next_work_cntr[3]), .B(next_work_cntr[2]), .C(
        next_work_cntr[1]), .D(\gt_357/A[0] ), .Y(n224) );
  NOR2BX2 U156 ( .AN(N141), .B(n220), .Y(next_work_cntr[3]) );
  AO22X2 U157 ( .A0(write_cntr[7]), .A1(n201), .B0(N273), .B1(n316), .Y(
        next_write_cntr[7]) );
  BUFX16 U158 ( .A(n614), .Y(cr_a[6]) );
  BUFX16 U159 ( .A(n601), .Y(im_a[9]) );
  NOR2X2 U160 ( .A(n220), .B(n332), .Y(next_work_cntr[8]) );
  NOR2BX2 U161 ( .AN(N153), .B(n221), .Y(next_work_cntr[15]) );
  NOR4X1 U162 ( .A(next_work_cntr[16]), .B(next_work_cntr[15]), .C(
        next_work_cntr[14]), .D(next_work_cntr[13]), .Y(n228) );
  AO22X2 U163 ( .A0(write_cntr[10]), .A1(n201), .B0(N276), .B1(n316), .Y(
        next_write_cntr[10]) );
  BUFX16 U164 ( .A(n615), .Y(cr_a[5]) );
  BUFX16 U165 ( .A(n602), .Y(im_a[8]) );
  NOR2X2 U166 ( .A(n220), .B(n333), .Y(next_work_cntr[5]) );
  NOR4X1 U167 ( .A(next_work_cntr[5]), .B(next_work_cntr[19]), .C(
        next_work_cntr[18]), .D(next_work_cntr[17]), .Y(n227) );
  NOR2BX2 U168 ( .AN(N149), .B(n221), .Y(next_work_cntr[11]) );
  NOR4X1 U169 ( .A(next_work_cntr[12]), .B(next_work_cntr[11]), .C(
        next_work_cntr[10]), .D(n225), .Y(n229) );
  AO22X2 U170 ( .A0(write_cntr[8]), .A1(n201), .B0(N274), .B1(n200), .Y(
        next_write_cntr[8]) );
  BUFX16 U171 ( .A(n616), .Y(cr_a[4]) );
  BUFX16 U172 ( .A(n603), .Y(im_a[7]) );
  NOR2X2 U173 ( .A(n220), .B(n331), .Y(next_work_cntr[9]) );
  NOR2BX2 U174 ( .AN(N154), .B(n221), .Y(next_work_cntr[16]) );
  AO22X2 U175 ( .A0(write_cntr[11]), .A1(n201), .B0(N277), .B1(n200), .Y(
        next_write_cntr[11]) );
  BUFX16 U176 ( .A(n612), .Y(cr_a[8]) );
  BUFX16 U177 ( .A(n604), .Y(im_a[6]) );
  NOR2BX2 U178 ( .AN(N150), .B(n221), .Y(next_work_cntr[12]) );
  NOR2BX2 U179 ( .AN(N144), .B(n220), .Y(next_work_cntr[6]) );
  AOI222X4 U180 ( .A0(n213), .A1(next_write_cntr[1]), .B0(write_addr[1]), .B1(
        n199), .C0(N720), .C1(n205), .Y(n272) );
  AO22X2 U181 ( .A0(write_cntr[6]), .A1(n201), .B0(N272), .B1(n200), .Y(
        next_write_cntr[6]) );
  BUFX16 U182 ( .A(n617), .Y(cr_a[3]) );
  BUFX16 U183 ( .A(n605), .Y(im_a[5]) );
  NOR3X2 U184 ( .A(n525), .B(state[2]), .C(n414), .Y(n545) );
  INVX1 U185 ( .A(state[0]), .Y(n414) );
  NOR4X2 U186 ( .A(n453), .B(init_time_mux_sel), .C(n432), .D(global_cntr[1]), 
        .Y(en_photo_num) );
  NOR2BX2 U187 ( .AN(N155), .B(n221), .Y(next_work_cntr[17]) );
  NOR2BX2 U188 ( .AN(N145), .B(n220), .Y(next_work_cntr[7]) );
  AOI222X4 U189 ( .A0(n213), .A1(n33), .B0(write_addr[2]), .B1(n199), .C0(N721), .C1(n205), .Y(n269) );
  AO22X2 U190 ( .A0(write_cntr[5]), .A1(n201), .B0(N271), .B1(n316), .Y(
        next_write_cntr[5]) );
  BUFX16 U191 ( .A(n618), .Y(cr_a[2]) );
  BUFX16 U192 ( .A(n606), .Y(im_a[4]) );
  NOR2BX2 U193 ( .AN(N151), .B(n221), .Y(next_work_cntr[13]) );
  NOR2BX2 U194 ( .AN(N156), .B(n220), .Y(next_work_cntr[18]) );
  NOR3X2 U195 ( .A(global_cntr[2]), .B(n454), .C(n432), .Y(N1425) );
  NOR3X2 U196 ( .A(state[0]), .B(state[2]), .C(n525), .Y(n503) );
  OAI222X1 U197 ( .A0(n198), .A1(n274), .B0(n307), .B1(n232), .C0(n308), .C1(
        n246), .Y(read_addr[0]) );
  AOI222X4 U198 ( .A0(n213), .A1(next_write_cntr[0]), .B0(write_addr[0]), .B1(
        n199), .C0(N719), .C1(n205), .Y(n308) );
  AO22X2 U199 ( .A0(write_cntr[3]), .A1(n201), .B0(N269), .B1(n316), .Y(
        next_write_cntr[3]) );
  BUFX16 U200 ( .A(n619), .Y(cr_a[1]) );
  BUFX16 U201 ( .A(n607), .Y(im_a[3]) );
  NOR2BX2 U202 ( .AN(N152), .B(n221), .Y(next_work_cntr[14]) );
  NOR2BX2 U203 ( .AN(N157), .B(n220), .Y(next_work_cntr[19]) );
  AO22X2 U204 ( .A0(write_cntr[1]), .A1(n201), .B0(N267), .B1(n316), .Y(
        next_write_cntr[1]) );
  NOR4X2 U205 ( .A(n455), .B(n453), .C(n434), .D(global_cntr[1]), .Y(N1447) );
  CLKINVX1 U206 ( .A(n537), .Y(next_state[0]) );
  OAI221XL U207 ( .A0(n573), .A1(n536), .B0(state[0]), .B1(n537), .C0(n538), 
        .Y(n325) );
  MXI2X2 U208 ( .A(n546), .B(n338), .S0(n503), .Y(n537) );
  AO22X2 U209 ( .A0(write_cntr[15]), .A1(n201), .B0(N281), .B1(n200), .Y(
        next_write_cntr[15]) );
  BUFX16 U210 ( .A(n620), .Y(cr_a[0]) );
  BUFX16 U211 ( .A(n609), .Y(im_a[1]) );
  NOR2BX2 U212 ( .AN(n428), .B(n419), .Y(n418) );
  NOR2BX2 U213 ( .AN(N138), .B(n220), .Y(\gt_357/A[0] ) );
  NOR2X2 U214 ( .A(n220), .B(n337), .Y(next_work_cntr[10]) );
  OAI21X1 U215 ( .A0(n551), .A1(n349), .B0(n552), .Y(n543) );
  AO22X2 U216 ( .A0(write_cntr[13]), .A1(n201), .B0(N279), .B1(n200), .Y(
        next_write_cntr[13]) );
  AO22X2 U217 ( .A0(write_cntr[16]), .A1(n201), .B0(N282), .B1(n316), .Y(
        next_write_cntr[16]) );
  AO22X4 U218 ( .A0(write_cntr[14]), .A1(n201), .B0(N280), .B1(n316), .Y(
        next_write_cntr[14]) );
  ADDHX1 U219 ( .A(s_1[3]), .B(\mult_236/n2 ), .CO(N640), .S(N639) );
  ADDHX1 U220 ( .A(m_1[3]), .B(\mult_234/n2 ), .CO(N604), .S(N603) );
  ADDHX1 U221 ( .A(h_1[3]), .B(\mult_232/n2 ), .CO(N568), .S(N567) );
  NOR4X2 U222 ( .A(init_time_mux_sel), .B(n433), .C(n434), .D(global_cntr[2]), 
        .Y(en_fb_addr) );
  OAI21X1 U223 ( .A0(n344), .A1(n345), .B0(n343), .Y(n342) );
  NOR3X4 U224 ( .A(n310), .B(read_cntr[0]), .C(n309), .Y(n278) );
  NAND2X2 U225 ( .A(n414), .B(en_so), .Y(n309) );
  OAI21X1 U226 ( .A0(next_state[1]), .A1(n573), .B0(next_state[0]), .Y(n324)
         );
  OAI221X4 U227 ( .A0(n544), .A1(n553), .B0(n13), .B1(n526), .C0(n17), .Y(n573) );
  OR2X2 U228 ( .A(next_en_si), .B(n221), .Y(_4_net_) );
  OAI22X1 U229 ( .A0(n339), .A1(n510), .B0(n329), .B1(n511), .Y(next_en_si) );
  BUFX16 U230 ( .A(n608), .Y(im_a[2]) );
  OA21X2 U231 ( .A0(n500), .A1(n212), .B0(n501), .Y(n611) );
  INVX16 U232 ( .A(n611), .Y(im_wen_n) );
  NAND2X2 U233 ( .A(n222), .B(im_wen_n), .Y(_6_net_) );
  INVX1 U234 ( .A(cr_x[1]), .Y(n494) );
  NAND2XL U235 ( .A(N657), .B(n149), .Y(n189) );
  NAND2XL U236 ( .A(N585), .B(n147), .Y(n193) );
  NAND2XL U237 ( .A(N621), .B(n148), .Y(n191) );
  NOR3XL U238 ( .A(N77), .B(N79), .C(N78), .Y(n508) );
  OR2XL U239 ( .A(next_work_cntr[3]), .B(\sub_358/carry[3] ), .Y(
        \sub_358/carry[4] ) );
  OR2XL U240 ( .A(next_work_cntr[1]), .B(\gt_357/A[0] ), .Y(\sub_358/carry[2] ) );
  OR2XL U241 ( .A(next_work_cntr[9]), .B(\sub_358/carry[9] ), .Y(
        \sub_358/carry[10] ) );
  OR2XL U242 ( .A(next_work_cntr[5]), .B(n146), .Y(\sub_358/carry[6] ) );
  OR2XL U243 ( .A(next_work_cntr[8]), .B(\sub_358/carry[8] ), .Y(
        \sub_358/carry[9] ) );
  OR2XL U244 ( .A(next_work_cntr[10]), .B(\sub_358/carry[10] ), .Y(
        \sub_358/carry[11] ) );
  OR2XL U245 ( .A(next_work_cntr[2]), .B(\sub_358/carry[2] ), .Y(
        \sub_358/carry[3] ) );
  AND2XL U246 ( .A(next_work_cntr[4]), .B(\sub_358/carry[4] ), .Y(n146) );
  NAND3XL U247 ( .A(cr_x[0]), .B(cr_x[1]), .C(n497), .Y(n491) );
  INVXL U248 ( .A(N24), .Y(n239) );
  INVX1 U249 ( .A(n542), .Y(next_state[1]) );
  MXI2XL U250 ( .A(n514), .B(n515), .S0(n238), .Y(n513) );
  OR2XL U251 ( .A(next_work_cntr[16]), .B(\sub_358/carry[16] ), .Y(
        \sub_358/carry[17] ) );
  OR2XL U252 ( .A(next_work_cntr[12]), .B(\sub_358/carry[12] ), .Y(
        \sub_358/carry[13] ) );
  OR2XL U253 ( .A(next_work_cntr[7]), .B(\sub_358/carry[7] ), .Y(
        \sub_358/carry[8] ) );
  OR2XL U254 ( .A(next_work_cntr[15]), .B(\sub_358/carry[15] ), .Y(
        \sub_358/carry[16] ) );
  OR2XL U255 ( .A(next_work_cntr[14]), .B(\sub_358/carry[14] ), .Y(
        \sub_358/carry[15] ) );
  OR2XL U256 ( .A(next_work_cntr[11]), .B(\sub_358/carry[11] ), .Y(
        \sub_358/carry[12] ) );
  OR2XL U257 ( .A(next_work_cntr[18]), .B(\sub_358/carry[18] ), .Y(
        \sub_358/carry[19] ) );
  OR2XL U258 ( .A(next_work_cntr[6]), .B(\sub_358/carry[6] ), .Y(
        \sub_358/carry[7] ) );
  OR2XL U259 ( .A(next_work_cntr[13]), .B(\sub_358/carry[13] ), .Y(
        \sub_358/carry[14] ) );
  OR2XL U260 ( .A(next_work_cntr[17]), .B(\sub_358/carry[17] ), .Y(
        \sub_358/carry[18] ) );
  OR4XL U261 ( .A(n239), .B(n240), .C(N22), .D(N23), .Y(n233) );
  NAND3XL U262 ( .A(n241), .B(n239), .C(N23), .Y(n235) );
  INVX1 U263 ( .A(n300), .Y(n232) );
  NAND2XL U264 ( .A(N567), .B(n153), .Y(n194) );
  NAND2XL U265 ( .A(N603), .B(n154), .Y(n192) );
  NAND2XL U266 ( .A(N639), .B(n155), .Y(n190) );
  NOR4XL U267 ( .A(next_work_cntr[9]), .B(next_work_cntr[8]), .C(
        next_work_cntr[7]), .D(next_work_cntr[6]), .Y(n226) );
  INVXL U268 ( .A(n240), .Y(n241) );
  INVXL U269 ( .A(n308), .Y(next_write_addr[0]) );
  INVXL U270 ( .A(n545), .Y(n553) );
  INVXL U271 ( .A(n272), .Y(next_write_addr[1]) );
  INVXL U272 ( .A(n266), .Y(next_write_addr[3]) );
  MXI2XL U273 ( .A(n212), .B(n502), .S0(n503), .Y(n501) );
  OAI211XL U274 ( .A0(n412), .A1(n504), .B0(n405), .C0(n328), .Y(n502) );
  INVXL U275 ( .A(n328), .Y(n338) );
  MXI2XL U276 ( .A(n305), .B(n306), .S0(n240), .Y(n304) );
  AOI21XL U277 ( .A0(N22), .A1(N23), .B0(N24), .Y(n305) );
  AOI21XL U278 ( .A0(N591), .A1(n461), .B0(n467), .Y(n475) );
  AOI21XL U279 ( .A0(N592), .A1(n461), .B0(n467), .Y(n472) );
  AOI21XL U280 ( .A0(N593), .A1(n461), .B0(n467), .Y(n469) );
  AOI21XL U281 ( .A0(N594), .A1(n461), .B0(n467), .Y(n465) );
  AOI22XL U282 ( .A0(N671), .A1(n460), .B0(N590), .B1(n461), .Y(n478) );
  AOI22XL U283 ( .A0(N569), .A1(n460), .B0(N569), .B1(n461), .Y(n487) );
  AOI22XL U284 ( .A0(N570), .A1(n460), .B0(N570), .B1(n461), .Y(n484) );
  AOI22XL U285 ( .A0(N571), .A1(n460), .B0(N571), .B1(n461), .Y(n481) );
  AOI22XL U286 ( .A0(N676), .A1(n460), .B0(N595), .B1(n461), .Y(n436) );
  AOI22XL U287 ( .A0(n418), .A1(n425), .B0(N77), .B1(n419), .Y(n424) );
  AOI22XL U288 ( .A0(n418), .A1(N390), .B0(N76), .B1(n419), .Y(n427) );
  AOI22XL U289 ( .A0(n418), .A1(n422), .B0(N78), .B1(n419), .Y(n421) );
  OAI211XL U290 ( .A0(n217), .A1(n417), .B0(n218), .C0(n418), .Y(n416) );
  NAND2XL U291 ( .A(N79), .B(n419), .Y(n415) );
  NAND4XL U292 ( .A(n535), .B(\gt_357/A[0] ), .C(n334), .D(n333), .Y(n533) );
  AOI22XL U293 ( .A0(write_addr[18]), .A1(n278), .B0(next_write_addr[18]), 
        .B1(n197), .Y(n281) );
  AOI2BB2XL U294 ( .B0(n261), .B1(next_write_addr[1]), .A0N(n271), .A1N(n195), 
        .Y(n270) );
  AOI2BB2XL U295 ( .B0(n261), .B1(next_write_addr[2]), .A0N(n268), .A1N(n195), 
        .Y(n267) );
  AOI2BB2XL U296 ( .B0(n261), .B1(next_write_addr[3]), .A0N(n265), .A1N(n195), 
        .Y(n264) );
  AOI2BB2XL U297 ( .B0(n261), .B1(next_write_addr[4]), .A0N(n262), .A1N(n195), 
        .Y(n260) );
  AOI22XL U298 ( .A0(n261), .A1(next_write_addr[13]), .B0(n289), .B1(
        write_addr[13]), .Y(n288) );
  AOI2BB2XL U299 ( .B0(write_addr[16]), .B1(n278), .A0N(n279), .A1N(n246), .Y(
        n287) );
  AOI22XL U300 ( .A0(n197), .A1(next_write_addr[13]), .B0(n278), .B1(
        write_addr[13]), .Y(n293) );
  AOI22XL U301 ( .A0(n261), .A1(next_write_addr[12]), .B0(n289), .B1(
        write_addr[12]), .Y(n290) );
  AOI2BB2XL U302 ( .B0(write_addr[17]), .B1(n278), .A0N(n275), .A1N(n246), .Y(
        n284) );
  AOI22XL U303 ( .A0(n197), .A1(next_write_addr[12]), .B0(n278), .B1(
        write_addr[12]), .Y(n296) );
  AOI22XL U304 ( .A0(write_addr[19]), .A1(n278), .B0(next_write_addr[19]), 
        .B1(n197), .Y(n277) );
  OAI2BB1XL U305 ( .A0N(n45), .A1N(n213), .B0(n313), .Y(next_write_addr[9]) );
  INVXL U306 ( .A(n257), .Y(next_write_addr[5]) );
  NAND3XL U307 ( .A(n525), .B(n536), .C(state[0]), .Y(n413) );
  AO22XL U308 ( .A0(next_write_cntr[18]), .A1(n213), .B0(n199), .B1(
        write_addr[18]), .Y(next_write_addr[18]) );
  AO22XL U309 ( .A0(n30), .A1(n213), .B0(n199), .B1(write_addr[19]), .Y(
        next_write_addr[19]) );
  MXI2XL U310 ( .A(n343), .B(n342), .S0(n379), .Y(next_photo[0]) );
  OR2XL U311 ( .A(n342), .B(n379), .Y(n341) );
  OA21XL U312 ( .A0(n328), .A1(n329), .B0(n330), .Y(n141) );
  XNOR2X1 U313 ( .A(work_cntr[17]), .B(\r898/carry[17] ), .Y(N1079) );
  AND4X1 U314 ( .A(n559), .B(n560), .C(n561), .D(n562), .Y(n142) );
  BUFX4 U315 ( .A(N1064), .Y(n217) );
  XNOR2X1 U316 ( .A(n74), .B(\sub_309/carry[18] ), .Y(N1045) );
  XNOR2X1 U317 ( .A(work_cntr[18]), .B(\r864/carry[18] ), .Y(N408) );
  XNOR2X1 U318 ( .A(n74), .B(\r902/carry[18] ), .Y(N1121) );
  AND2X2 U319 ( .A(N698), .B(n144), .Y(n143) );
  AND2X2 U320 ( .A(N697), .B(n145), .Y(n144) );
  INVX3 U321 ( .A(n490), .Y(n462) );
  AND2X2 U322 ( .A(N696), .B(\add_0_root_add_0_root_add_269_2/carry[4] ), .Y(
        n145) );
  CLKBUFX3 U323 ( .A(n458), .Y(n211) );
  NOR3BXL U324 ( .AN(n493), .B(n494), .C(n495), .Y(n458) );
  INVX3 U325 ( .A(n491), .Y(n463) );
  INVX3 U326 ( .A(n489), .Y(n461) );
  XOR2XL U327 ( .A(N585), .B(n147), .Y(N594) );
  XOR2XL U328 ( .A(N657), .B(n149), .Y(N666) );
  XOR2XL U329 ( .A(N621), .B(n148), .Y(N630) );
  XNOR2X1 U330 ( .A(N586), .B(n193), .Y(N595) );
  XNOR2X1 U331 ( .A(N658), .B(n189), .Y(N667) );
  XNOR2X1 U332 ( .A(N622), .B(n191), .Y(N631) );
  CLKBUFX3 U333 ( .A(n459), .Y(n209) );
  NOR3BXL U334 ( .AN(n493), .B(cr_x[0]), .C(cr_x[1]), .Y(n459) );
  CLKBUFX3 U335 ( .A(n457), .Y(n210) );
  NOR3BXL U336 ( .AN(n493), .B(cr_x[0]), .C(n494), .Y(n457) );
  XNOR2X1 U337 ( .A(next_work_cntr[10]), .B(\sub_358/carry[10] ), .Y(N1210) );
  XNOR2X1 U338 ( .A(next_work_cntr[9]), .B(\sub_358/carry[9] ), .Y(N1209) );
  XNOR2X1 U339 ( .A(next_work_cntr[8]), .B(\sub_358/carry[8] ), .Y(N1208) );
  XNOR2X1 U340 ( .A(next_work_cntr[5]), .B(n146), .Y(N1205) );
  XOR2X1 U341 ( .A(next_work_cntr[4]), .B(\sub_358/carry[4] ), .Y(N1204) );
  XNOR2X1 U342 ( .A(next_work_cntr[3]), .B(\sub_358/carry[3] ), .Y(N1203) );
  AND2X2 U343 ( .A(N584), .B(n156), .Y(n147) );
  AND2X2 U344 ( .A(N620), .B(n157), .Y(n148) );
  AND2X2 U345 ( .A(N656), .B(n158), .Y(n149) );
  XOR2X1 U346 ( .A(N565), .B(\add_232/carry[5] ), .Y(N574) );
  XOR2X1 U347 ( .A(N601), .B(\add_234/carry[5] ), .Y(N610) );
  XOR2X1 U348 ( .A(N584), .B(n156), .Y(N593) );
  XOR2X1 U349 ( .A(N656), .B(n158), .Y(N665) );
  XOR2X1 U350 ( .A(N637), .B(\add_236/carry[5] ), .Y(N646) );
  XOR2X1 U351 ( .A(N620), .B(n157), .Y(N629) );
  AND2X2 U352 ( .A(N565), .B(\add_232/carry[5] ), .Y(n150) );
  AND2X2 U353 ( .A(N601), .B(\add_234/carry[5] ), .Y(n151) );
  AND2X2 U354 ( .A(N637), .B(\add_236/carry[5] ), .Y(n152) );
  XNOR2X1 U355 ( .A(next_work_cntr[2]), .B(\sub_358/carry[2] ), .Y(N1202) );
  XNOR2X1 U356 ( .A(next_work_cntr[1]), .B(\gt_357/A[0] ), .Y(N1201) );
  BUFX4 U357 ( .A(n326), .Y(n202) );
  NOR2X1 U358 ( .A(n329), .B(n338), .Y(n326) );
  OR2X2 U359 ( .A(n202), .B(n204), .Y(n316) );
  BUFX4 U360 ( .A(n312), .Y(n213) );
  NOR2XL U361 ( .A(next_state[0]), .B(n542), .Y(n312) );
  CLKBUFX3 U362 ( .A(n314), .Y(n205) );
  NOR2XL U363 ( .A(n324), .B(n221), .Y(n314) );
  OR2X2 U364 ( .A(n202), .B(n204), .Y(n200) );
  XNOR2X1 U365 ( .A(next_work_cntr[17]), .B(\sub_358/carry[17] ), .Y(N1217) );
  XNOR2X1 U366 ( .A(next_work_cntr[18]), .B(\sub_358/carry[18] ), .Y(N1218) );
  XNOR2X1 U367 ( .A(next_work_cntr[19]), .B(\sub_358/carry[19] ), .Y(N1219) );
  XNOR2X1 U368 ( .A(next_work_cntr[16]), .B(\sub_358/carry[16] ), .Y(N1216) );
  XNOR2X1 U369 ( .A(next_work_cntr[15]), .B(\sub_358/carry[15] ), .Y(N1215) );
  XNOR2X1 U370 ( .A(next_work_cntr[14]), .B(\sub_358/carry[14] ), .Y(N1214) );
  CLKBUFX3 U371 ( .A(n248), .Y(n196) );
  NAND2XL U372 ( .A(n302), .B(n300), .Y(n248) );
  CLKBUFX3 U373 ( .A(n250), .Y(n195) );
  NAND2XL U374 ( .A(n300), .B(n301), .Y(n250) );
  XNOR2X1 U375 ( .A(next_work_cntr[13]), .B(\sub_358/carry[13] ), .Y(N1213) );
  XNOR2X1 U376 ( .A(next_work_cntr[12]), .B(\sub_358/carry[12] ), .Y(N1212) );
  BUFX4 U377 ( .A(n364), .Y(n206) );
  OAI21XL U378 ( .A0(n309), .A1(n405), .B0(n406), .Y(n364) );
  XNOR2X1 U379 ( .A(next_work_cntr[11]), .B(\sub_358/carry[11] ), .Y(N1211) );
  BUFX4 U380 ( .A(n363), .Y(n207) );
  OAI21XL U381 ( .A0(n238), .A1(n231), .B0(n409), .Y(n363) );
  XNOR2X1 U382 ( .A(next_work_cntr[7]), .B(\sub_358/carry[7] ), .Y(N1207) );
  XNOR2X1 U383 ( .A(next_work_cntr[6]), .B(\sub_358/carry[6] ), .Y(N1206) );
  BUFX4 U384 ( .A(n315), .Y(n199) );
  NOR3BXL U385 ( .AN(n324), .B(n213), .C(n221), .Y(n315) );
  XOR2XL U386 ( .A(N567), .B(n153), .Y(N576) );
  XOR2XL U387 ( .A(N603), .B(n154), .Y(N612) );
  XOR2XL U388 ( .A(N639), .B(n155), .Y(N648) );
  XNOR2X1 U389 ( .A(N568), .B(n194), .Y(N577) );
  XNOR2X1 U390 ( .A(N604), .B(n192), .Y(N613) );
  AND2X2 U391 ( .A(N566), .B(n150), .Y(n153) );
  AND2X2 U392 ( .A(N602), .B(n151), .Y(n154) );
  AND2X2 U393 ( .A(N638), .B(n152), .Y(n155) );
  AND2X2 U394 ( .A(N583), .B(\add_233/carry[5] ), .Y(n156) );
  AND2X2 U395 ( .A(N619), .B(\add_235/carry[5] ), .Y(n157) );
  XNOR2X1 U396 ( .A(N640), .B(n190), .Y(N649) );
  XOR2X1 U397 ( .A(N566), .B(n150), .Y(N575) );
  XOR2X1 U398 ( .A(N602), .B(n151), .Y(N611) );
  XOR2X1 U399 ( .A(N583), .B(\add_233/carry[5] ), .Y(N592) );
  XOR2X1 U400 ( .A(N655), .B(\add_237/carry[5] ), .Y(N664) );
  XOR2X1 U401 ( .A(N638), .B(n152), .Y(N647) );
  XOR2X1 U402 ( .A(N619), .B(\add_235/carry[5] ), .Y(N628) );
  AND2X2 U403 ( .A(N655), .B(\add_237/carry[5] ), .Y(n158) );
  XOR2X1 U404 ( .A(N671), .B(N563), .Y(N572) );
  XOR2X1 U405 ( .A(N671), .B(N599), .Y(N608) );
  XOR2X1 U406 ( .A(N671), .B(N635), .Y(N644) );
  INVX3 U407 ( .A(n197), .Y(n246) );
  NAND2X2 U408 ( .A(n330), .B(n329), .Y(n352) );
  INVX4 U409 ( .A(n141), .Y(n201) );
  INVX3 U410 ( .A(n222), .Y(n221) );
  CLKBUFX3 U411 ( .A(n327), .Y(n204) );
  NOR2BX1 U412 ( .AN(n205), .B(n353), .Y(n327) );
  BUFX4 U413 ( .A(n362), .Y(n214) );
  CLKINVX1 U414 ( .A(n413), .Y(n362) );
  OR2X1 U415 ( .A(n218), .B(n159), .Y(\sub_309/carry[4] ) );
  AND2X2 U416 ( .A(n217), .B(n160), .Y(n159) );
  AND2X2 U417 ( .A(n216), .B(n219), .Y(n160) );
  INVX3 U418 ( .A(n222), .Y(n220) );
  OR2X1 U419 ( .A(n218), .B(n161), .Y(\r864/carry[4] ) );
  AND2X2 U420 ( .A(n217), .B(n162), .Y(n161) );
  AND2X2 U421 ( .A(n216), .B(n219), .Y(n162) );
  XNOR2X1 U422 ( .A(n218), .B(n159), .Y(N1030) );
  OR2X1 U423 ( .A(n218), .B(n163), .Y(\r902/carry[4] ) );
  AND2X2 U424 ( .A(n217), .B(n216), .Y(n163) );
  XOR2X1 U425 ( .A(n217), .B(n160), .Y(N1029) );
  XOR2X1 U426 ( .A(n216), .B(n219), .Y(N1028) );
  XNOR2X1 U427 ( .A(n218), .B(n161), .Y(N393) );
  XOR2X1 U428 ( .A(N671), .B(N581), .Y(N590) );
  XOR2X1 U429 ( .A(N671), .B(N617), .Y(N626) );
  XOR2X1 U430 ( .A(n217), .B(n162), .Y(N392) );
  XOR2X1 U431 ( .A(N671), .B(N653), .Y(N662) );
  CLKBUFX3 U432 ( .A(n243), .Y(n198) );
  INVXL U433 ( .A(n278), .Y(n243) );
  XOR2X1 U434 ( .A(n216), .B(n219), .Y(N391) );
  CLKBUFX3 U435 ( .A(n252), .Y(n197) );
  NOR3XL U436 ( .A(n309), .B(n310), .C(n311), .Y(n252) );
  BUFX4 U437 ( .A(n359), .Y(n208) );
  NAND3XL U438 ( .A(n309), .B(n212), .C(n413), .Y(n359) );
  XNOR2X1 U439 ( .A(N811), .B(n188), .Y(N993) );
  NAND2X1 U440 ( .A(N810), .B(n165), .Y(n188) );
  AND2X2 U441 ( .A(N808), .B(\add_0_root_add_296_2/carry[16] ), .Y(n164) );
  AND2X2 U442 ( .A(N809), .B(n164), .Y(n165) );
  XNOR2X1 U443 ( .A(N806), .B(\add_0_root_add_296_2/carry[14] ), .Y(N988) );
  XNOR2X1 U444 ( .A(N807), .B(\add_0_root_add_296_2/carry[15] ), .Y(N989) );
  XOR2X1 U445 ( .A(N808), .B(\add_0_root_add_296_2/carry[16] ), .Y(N990) );
  XOR2X1 U446 ( .A(N809), .B(n164), .Y(N991) );
  XOR2X1 U447 ( .A(N810), .B(n165), .Y(N992) );
  XNOR2X1 U448 ( .A(n218), .B(n163), .Y(N1106) );
  OR2X1 U449 ( .A(N805), .B(n166), .Y(\add_0_root_add_296_2/carry[14] ) );
  OR2X1 U450 ( .A(N806), .B(\add_0_root_add_296_2/carry[14] ), .Y(
        \add_0_root_add_296_2/carry[15] ) );
  OR2X1 U451 ( .A(N796), .B(N795), .Y(\add_0_root_add_296_2/carry[5] ) );
  OR2X1 U452 ( .A(N799), .B(n167), .Y(\add_0_root_add_296_2/carry[8] ) );
  OR2X1 U453 ( .A(N803), .B(n168), .Y(\add_0_root_add_296_2/carry[12] ) );
  BUFX4 U454 ( .A(n621), .Y(si_sel) );
  AND2X2 U455 ( .A(N804), .B(\add_0_root_add_296_2/carry[12] ), .Y(n166) );
  AND2X2 U456 ( .A(N798), .B(n169), .Y(n167) );
  AND2X2 U457 ( .A(N802), .B(n171), .Y(n168) );
  AND2X2 U458 ( .A(N797), .B(\add_0_root_add_296_2/carry[5] ), .Y(n169) );
  AND2X2 U459 ( .A(N800), .B(\add_0_root_add_296_2/carry[8] ), .Y(n170) );
  AND2X2 U460 ( .A(N801), .B(n170), .Y(n171) );
  OR2X1 U461 ( .A(N807), .B(\add_0_root_add_296_2/carry[15] ), .Y(
        \add_0_root_add_296_2/carry[16] ) );
  XOR2X1 U462 ( .A(N804), .B(\add_0_root_add_296_2/carry[12] ), .Y(N986) );
  XNOR2X1 U463 ( .A(N803), .B(n168), .Y(N985) );
  XNOR2X1 U464 ( .A(N805), .B(n166), .Y(N987) );
  XOR2X1 U465 ( .A(N801), .B(n170), .Y(N983) );
  XOR2X1 U466 ( .A(N802), .B(n171), .Y(N984) );
  INVX4 U467 ( .A(n18), .Y(n203) );
  XOR2X1 U468 ( .A(n217), .B(n216), .Y(N1105) );
  XNOR2X1 U469 ( .A(N796), .B(N795), .Y(N978) );
  XOR2X1 U470 ( .A(N797), .B(\add_0_root_add_296_2/carry[5] ), .Y(N979) );
  XOR2X1 U471 ( .A(N800), .B(\add_0_root_add_296_2/carry[8] ), .Y(N982) );
  XNOR2X1 U472 ( .A(N799), .B(n167), .Y(N981) );
  XOR2X1 U473 ( .A(N798), .B(n169), .Y(N980) );
  CLKINVX1 U474 ( .A(N795), .Y(N977) );
  CLKINVX1 U475 ( .A(n216), .Y(N1104) );
  XNOR2X1 U476 ( .A(n74), .B(\r898/carry[18] ), .Y(N1080) );
  XNOR2X1 U477 ( .A(n85), .B(\r898/carry[19] ), .Y(N1081) );
  OR2X1 U478 ( .A(n96), .B(\r898/carry[6] ), .Y(\r898/carry[7] ) );
  OR2X1 U479 ( .A(n100), .B(\r898/carry[7] ), .Y(\r898/carry[8] ) );
  OR2X1 U480 ( .A(n98), .B(\r898/carry[8] ), .Y(\r898/carry[9] ) );
  OR2X1 U481 ( .A(n102), .B(\r898/carry[9] ), .Y(\r898/carry[10] ) );
  OR2X1 U482 ( .A(n77), .B(\r898/carry[10] ), .Y(\r898/carry[11] ) );
  OR2X1 U483 ( .A(n87), .B(\r898/carry[11] ), .Y(\r898/carry[12] ) );
  OR2X1 U484 ( .A(n92), .B(\r898/carry[12] ), .Y(\r898/carry[13] ) );
  OR2X1 U485 ( .A(n81), .B(\r898/carry[13] ), .Y(\r898/carry[14] ) );
  OR2X1 U486 ( .A(n90), .B(\r898/carry[14] ), .Y(\r898/carry[15] ) );
  OR2X1 U487 ( .A(n94), .B(\r898/carry[15] ), .Y(\r898/carry[16] ) );
  OR2X1 U488 ( .A(n79), .B(\r898/carry[16] ), .Y(\r898/carry[17] ) );
  OR2X1 U489 ( .A(work_cntr[17]), .B(\r898/carry[17] ), .Y(\r898/carry[18] )
         );
  OR2X1 U490 ( .A(n74), .B(\r898/carry[18] ), .Y(\r898/carry[19] ) );
  XNOR2X1 U491 ( .A(n79), .B(\r898/carry[16] ), .Y(N1078) );
  XNOR2X1 U492 ( .A(n94), .B(\r898/carry[15] ), .Y(N1077) );
  XNOR2X1 U493 ( .A(n90), .B(\r898/carry[14] ), .Y(N1076) );
  XNOR2X1 U494 ( .A(n81), .B(\r898/carry[13] ), .Y(N1075) );
  XOR2X1 U495 ( .A(global_cntr[18]), .B(n186), .Y(N1012) );
  XOR2X1 U496 ( .A(global_cntr[19]), .B(n187), .Y(N1013) );
  CLKINVX1 U497 ( .A(n325), .Y(n222) );
  XOR2X1 U498 ( .A(global_cntr[13]), .B(n181), .Y(N1007) );
  XOR2X1 U499 ( .A(global_cntr[15]), .B(n183), .Y(N1009) );
  XOR2X1 U500 ( .A(global_cntr[16]), .B(n184), .Y(N1010) );
  XOR2X1 U501 ( .A(global_cntr[14]), .B(n182), .Y(N1008) );
  XOR2X1 U502 ( .A(global_cntr[17]), .B(n185), .Y(N1011) );
  XNOR2X1 U503 ( .A(work_cntr[12]), .B(\r898/carry[12] ), .Y(N1074) );
  XOR2X1 U504 ( .A(global_cntr[8]), .B(n176), .Y(N1002) );
  XOR2X1 U505 ( .A(global_cntr[12]), .B(n180), .Y(N1006) );
  XOR2X1 U506 ( .A(N697), .B(n145), .Y(N724) );
  XOR2X1 U507 ( .A(N692), .B(\add_0_root_add_0_root_add_269_2/A[0] ), .Y(N719)
         );
  XOR2X1 U508 ( .A(N696), .B(\add_0_root_add_0_root_add_269_2/carry[4] ), .Y(
        N723) );
  XOR2X1 U509 ( .A(N698), .B(n144), .Y(N725) );
  XOR2X1 U510 ( .A(N699), .B(n143), .Y(N726) );
  XOR2X1 U511 ( .A(global_cntr[9]), .B(n177), .Y(N1003) );
  XOR2X1 U512 ( .A(global_cntr[10]), .B(n178), .Y(N1004) );
  XOR2X1 U513 ( .A(global_cntr[11]), .B(n179), .Y(N1005) );
  INVX4 U514 ( .A(n142), .Y(n215) );
  XNOR2X1 U515 ( .A(n87), .B(\r898/carry[11] ), .Y(N1073) );
  XOR2X1 U516 ( .A(global_cntr[6]), .B(n174), .Y(N1000) );
  XOR2X1 U517 ( .A(global_cntr[7]), .B(n175), .Y(N1001) );
  XOR2X1 U518 ( .A(global_cntr[3]), .B(\add_298/carry[3] ), .Y(N997) );
  XOR2X1 U519 ( .A(global_cntr[4]), .B(n172), .Y(N998) );
  XOR2X1 U520 ( .A(global_cntr[5]), .B(n173), .Y(N999) );
  XNOR2X1 U521 ( .A(n77), .B(\r898/carry[10] ), .Y(N1072) );
  XNOR2X1 U522 ( .A(n85), .B(\sub_309/carry[19] ), .Y(N1046) );
  OR2X1 U523 ( .A(work_cntr[4]), .B(\sub_309/carry[4] ), .Y(\sub_309/carry[5] ) );
  OR2X1 U524 ( .A(n83), .B(\sub_309/carry[5] ), .Y(\sub_309/carry[6] ) );
  OR2X1 U525 ( .A(n96), .B(\sub_309/carry[6] ), .Y(\sub_309/carry[7] ) );
  OR2X1 U526 ( .A(n100), .B(\sub_309/carry[7] ), .Y(\sub_309/carry[8] ) );
  OR2X1 U527 ( .A(n98), .B(\sub_309/carry[8] ), .Y(\sub_309/carry[9] ) );
  OR2X1 U528 ( .A(n102), .B(\sub_309/carry[9] ), .Y(\sub_309/carry[10] ) );
  OR2X1 U529 ( .A(n77), .B(\sub_309/carry[10] ), .Y(\sub_309/carry[11] ) );
  OR2X1 U530 ( .A(n87), .B(\sub_309/carry[11] ), .Y(\sub_309/carry[12] ) );
  OR2X1 U531 ( .A(n92), .B(\sub_309/carry[12] ), .Y(\sub_309/carry[13] ) );
  OR2X1 U532 ( .A(n81), .B(\sub_309/carry[13] ), .Y(\sub_309/carry[14] ) );
  OR2X1 U533 ( .A(n90), .B(\sub_309/carry[14] ), .Y(\sub_309/carry[15] ) );
  OR2X1 U534 ( .A(n94), .B(\sub_309/carry[15] ), .Y(\sub_309/carry[16] ) );
  OR2X1 U535 ( .A(n79), .B(\sub_309/carry[16] ), .Y(\sub_309/carry[17] ) );
  OR2X1 U536 ( .A(work_cntr[17]), .B(\sub_309/carry[17] ), .Y(
        \sub_309/carry[18] ) );
  OR2X1 U537 ( .A(n74), .B(\sub_309/carry[18] ), .Y(\sub_309/carry[19] ) );
  BUFX4 U538 ( .A(N1062), .Y(n219) );
  BUFX4 U539 ( .A(N1063), .Y(n216) );
  BUFX4 U540 ( .A(N1065), .Y(n218) );
  XOR2X1 U541 ( .A(curr_photo[0]), .B(global_cntr[1]), .Y(N995) );
  XNOR2X1 U542 ( .A(work_cntr[17]), .B(\sub_309/carry[17] ), .Y(N1044) );
  XNOR2X1 U543 ( .A(n79), .B(\sub_309/carry[16] ), .Y(N1043) );
  XNOR2X1 U544 ( .A(n102), .B(\r898/carry[9] ), .Y(N1071) );
  XNOR2X1 U545 ( .A(n94), .B(\sub_309/carry[15] ), .Y(N1042) );
  XNOR2X1 U546 ( .A(n98), .B(\r898/carry[8] ), .Y(N1070) );
  XNOR2X1 U547 ( .A(work_cntr[14]), .B(\sub_309/carry[14] ), .Y(N1041) );
  XNOR2X1 U548 ( .A(n100), .B(\r898/carry[7] ), .Y(N1069) );
  XNOR2X1 U549 ( .A(work_cntr[13]), .B(\sub_309/carry[13] ), .Y(N1040) );
  XNOR2X1 U550 ( .A(n92), .B(\sub_309/carry[12] ), .Y(N1039) );
  XNOR2X1 U551 ( .A(n96), .B(\r898/carry[6] ), .Y(N1068) );
  XNOR2X1 U552 ( .A(n83), .B(work_cntr[4]), .Y(N1067) );
  XNOR2X1 U553 ( .A(n88), .B(\sub_309/carry[11] ), .Y(N1038) );
  CLKINVX1 U554 ( .A(work_cntr[4]), .Y(N1066) );
  XNOR2X1 U555 ( .A(n76), .B(\sub_309/carry[10] ), .Y(N1037) );
  XNOR2X1 U556 ( .A(n102), .B(\sub_309/carry[9] ), .Y(N1036) );
  XNOR2X1 U557 ( .A(work_cntr[19]), .B(\r864/carry[19] ), .Y(N409) );
  OR2X1 U558 ( .A(work_cntr[4]), .B(\r864/carry[4] ), .Y(\r864/carry[5] ) );
  OR2X1 U559 ( .A(work_cntr[5]), .B(\r864/carry[5] ), .Y(\r864/carry[6] ) );
  OR2X1 U560 ( .A(work_cntr[6]), .B(\r864/carry[6] ), .Y(\r864/carry[7] ) );
  OR2X1 U561 ( .A(work_cntr[7]), .B(\r864/carry[7] ), .Y(\r864/carry[8] ) );
  OR2X1 U562 ( .A(work_cntr[8]), .B(\r864/carry[8] ), .Y(\r864/carry[9] ) );
  OR2X1 U563 ( .A(work_cntr[9]), .B(\r864/carry[9] ), .Y(\r864/carry[10] ) );
  OR2X1 U564 ( .A(work_cntr[10]), .B(\r864/carry[10] ), .Y(\r864/carry[11] )
         );
  OR2X1 U565 ( .A(work_cntr[11]), .B(\r864/carry[11] ), .Y(\r864/carry[12] )
         );
  OR2X1 U566 ( .A(work_cntr[12]), .B(\r864/carry[12] ), .Y(\r864/carry[13] )
         );
  OR2X1 U567 ( .A(work_cntr[13]), .B(\r864/carry[13] ), .Y(\r864/carry[14] )
         );
  OR2X1 U568 ( .A(work_cntr[14]), .B(\r864/carry[14] ), .Y(\r864/carry[15] )
         );
  OR2X1 U569 ( .A(work_cntr[15]), .B(\r864/carry[15] ), .Y(\r864/carry[16] )
         );
  OR2X1 U570 ( .A(work_cntr[16]), .B(\r864/carry[16] ), .Y(\r864/carry[17] )
         );
  OR2X1 U571 ( .A(work_cntr[17]), .B(\r864/carry[17] ), .Y(\r864/carry[18] )
         );
  OR2X1 U572 ( .A(work_cntr[18]), .B(\r864/carry[18] ), .Y(\r864/carry[19] )
         );
  XNOR2X1 U573 ( .A(work_cntr[17]), .B(\r864/carry[17] ), .Y(N407) );
  XNOR2X1 U574 ( .A(n98), .B(\sub_309/carry[8] ), .Y(N1035) );
  XNOR2X1 U575 ( .A(work_cntr[16]), .B(\r864/carry[16] ), .Y(N406) );
  XNOR2X1 U576 ( .A(n100), .B(\sub_309/carry[7] ), .Y(N1034) );
  XNOR2X1 U577 ( .A(n94), .B(\r864/carry[15] ), .Y(N405) );
  XNOR2X1 U578 ( .A(n96), .B(\sub_309/carry[6] ), .Y(N1033) );
  BUFX4 U579 ( .A(n234), .Y(n212) );
  NAND2XL U580 ( .A(state[0]), .B(en_so), .Y(n234) );
  XNOR2X1 U581 ( .A(work_cntr[14]), .B(\r864/carry[14] ), .Y(N404) );
  XNOR2X1 U582 ( .A(n83), .B(\sub_309/carry[5] ), .Y(N1032) );
  XNOR2X1 U583 ( .A(n81), .B(\r864/carry[13] ), .Y(N403) );
  XNOR2X1 U584 ( .A(work_cntr[4]), .B(\sub_309/carry[4] ), .Y(N1031) );
  XNOR2X1 U585 ( .A(work_cntr[12]), .B(\r864/carry[12] ), .Y(N402) );
  XNOR2X1 U586 ( .A(work_cntr[11]), .B(\r864/carry[11] ), .Y(N401) );
  XNOR2X1 U587 ( .A(n85), .B(\r902/carry[19] ), .Y(N1122) );
  OR2X1 U588 ( .A(work_cntr[4]), .B(\r902/carry[4] ), .Y(\r902/carry[5] ) );
  OR2X1 U589 ( .A(n83), .B(\r902/carry[5] ), .Y(\r902/carry[6] ) );
  OR2X1 U590 ( .A(n96), .B(\r902/carry[6] ), .Y(\r902/carry[7] ) );
  OR2X1 U591 ( .A(n100), .B(\r902/carry[7] ), .Y(\r902/carry[8] ) );
  OR2X1 U592 ( .A(n98), .B(\r902/carry[8] ), .Y(\r902/carry[9] ) );
  OR2X1 U593 ( .A(n102), .B(\r902/carry[9] ), .Y(\r902/carry[10] ) );
  OR2X1 U594 ( .A(n77), .B(\r902/carry[10] ), .Y(\r902/carry[11] ) );
  OR2X1 U595 ( .A(n87), .B(\r902/carry[11] ), .Y(\r902/carry[12] ) );
  OR2X1 U596 ( .A(n92), .B(\r902/carry[12] ), .Y(\r902/carry[13] ) );
  OR2X1 U597 ( .A(work_cntr[13]), .B(\r902/carry[13] ), .Y(\r902/carry[14] )
         );
  OR2X1 U598 ( .A(n90), .B(\r902/carry[14] ), .Y(\r902/carry[15] ) );
  OR2X1 U599 ( .A(work_cntr[15]), .B(\r902/carry[15] ), .Y(\r902/carry[16] )
         );
  OR2X1 U600 ( .A(n79), .B(\r902/carry[16] ), .Y(\r902/carry[17] ) );
  OR2X1 U601 ( .A(work_cntr[17]), .B(\r902/carry[17] ), .Y(\r902/carry[18] )
         );
  OR2X1 U602 ( .A(n74), .B(\r902/carry[18] ), .Y(\r902/carry[19] ) );
  XNOR2X1 U603 ( .A(work_cntr[17]), .B(\r902/carry[17] ), .Y(N1120) );
  XNOR2X1 U604 ( .A(work_cntr[16]), .B(\r902/carry[16] ), .Y(N1119) );
  XNOR2X1 U605 ( .A(work_cntr[10]), .B(\r864/carry[10] ), .Y(N400) );
  XNOR2X1 U606 ( .A(work_cntr[15]), .B(\r902/carry[15] ), .Y(N1118) );
  XNOR2X1 U607 ( .A(n102), .B(\r864/carry[9] ), .Y(N399) );
  XNOR2X1 U608 ( .A(n98), .B(\r864/carry[8] ), .Y(N398) );
  XNOR2X1 U609 ( .A(n90), .B(\r902/carry[14] ), .Y(N1117) );
  XNOR2X1 U610 ( .A(n81), .B(\r902/carry[13] ), .Y(N1116) );
  XNOR2X1 U611 ( .A(n100), .B(\r864/carry[7] ), .Y(N397) );
  XNOR2X1 U612 ( .A(n96), .B(\r864/carry[6] ), .Y(N396) );
  XNOR2X1 U613 ( .A(work_cntr[12]), .B(\r902/carry[12] ), .Y(N1115) );
  XNOR2X1 U614 ( .A(n87), .B(\r902/carry[11] ), .Y(N1114) );
  XNOR2X1 U615 ( .A(n83), .B(\r864/carry[5] ), .Y(N395) );
  XNOR2X1 U616 ( .A(work_cntr[4]), .B(\r864/carry[4] ), .Y(N394) );
  XNOR2X1 U617 ( .A(n77), .B(\r902/carry[10] ), .Y(N1113) );
  XNOR2X1 U618 ( .A(n102), .B(\r902/carry[9] ), .Y(N1112) );
  XNOR2X1 U619 ( .A(n98), .B(\r902/carry[8] ), .Y(N1111) );
  XNOR2X1 U620 ( .A(n100), .B(\r902/carry[7] ), .Y(N1110) );
  XNOR2X1 U621 ( .A(n96), .B(\r902/carry[6] ), .Y(N1109) );
  XNOR2X1 U622 ( .A(n83), .B(\r902/carry[5] ), .Y(N1108) );
  XNOR2X1 U623 ( .A(work_cntr[4]), .B(\r902/carry[4] ), .Y(N1107) );
  AND2X2 U624 ( .A(global_cntr[3]), .B(\add_298/carry[3] ), .Y(n172) );
  AND2X2 U625 ( .A(global_cntr[4]), .B(n172), .Y(n173) );
  AND2X2 U626 ( .A(global_cntr[5]), .B(n173), .Y(n174) );
  AND2X2 U627 ( .A(global_cntr[6]), .B(n174), .Y(n175) );
  AND2X2 U628 ( .A(global_cntr[7]), .B(n175), .Y(n176) );
  AND2X2 U629 ( .A(global_cntr[8]), .B(n176), .Y(n177) );
  AND2X2 U630 ( .A(global_cntr[9]), .B(n177), .Y(n178) );
  AND2X2 U631 ( .A(global_cntr[10]), .B(n178), .Y(n179) );
  AND2X2 U632 ( .A(global_cntr[11]), .B(n179), .Y(n180) );
  AND2X2 U633 ( .A(global_cntr[12]), .B(n180), .Y(n181) );
  AND2X2 U634 ( .A(global_cntr[13]), .B(n181), .Y(n182) );
  AND2X2 U635 ( .A(global_cntr[14]), .B(n182), .Y(n183) );
  AND2X2 U636 ( .A(global_cntr[15]), .B(n183), .Y(n184) );
  AND2X2 U637 ( .A(global_cntr[16]), .B(n184), .Y(n185) );
  AND2X2 U638 ( .A(global_cntr[17]), .B(n185), .Y(n186) );
  AND2X2 U639 ( .A(global_cntr[18]), .B(n186), .Y(n187) );
  CLKINVX1 U640 ( .A(\gt_357/A[0] ), .Y(N1200) );
  CLKINVX1 U641 ( .A(n219), .Y(N390) );
  NOR2BX1 U642 ( .AN(next_work_cntr[4]), .B(n224), .Y(n225) );
  NAND4X1 U643 ( .A(n229), .B(n228), .C(n227), .D(n226), .Y(N1198) );
  AOI31X1 U644 ( .A0(n235), .A1(n233), .A2(n236), .B0(n232), .Y(so_mux_sel[0])
         );
  NAND2BX1 U645 ( .AN(n237), .B(n238), .Y(n236) );
  OAI222XL U646 ( .A0(n232), .A1(n242), .B0(n198), .B1(n244), .C0(n245), .C1(
        n246), .Y(read_addr[9]) );
  OAI221XL U647 ( .A0(n247), .A1(n196), .B0(n249), .B1(n195), .C0(n251), .Y(
        read_addr[8]) );
  AOI2BB2X1 U648 ( .B0(n197), .B1(next_write_addr[8]), .A0N(n198), .A1N(n253), 
        .Y(n251) );
  CLKINVX1 U649 ( .A(next_write_addr[7]), .Y(n247) );
  OAI221XL U650 ( .A0(n254), .A1(n196), .B0(n195), .B1(n255), .C0(n256), .Y(
        read_addr[7]) );
  AOI2BB2X1 U651 ( .B0(n197), .B1(next_write_addr[7]), .A0N(n198), .A1N(n249), 
        .Y(n256) );
  CLKINVX1 U652 ( .A(write_addr[7]), .Y(n249) );
  CLKINVX1 U653 ( .A(next_write_addr[6]), .Y(n254) );
  OAI221XL U654 ( .A0(n257), .A1(n196), .B0(n195), .B1(n258), .C0(n259), .Y(
        read_addr[6]) );
  AOI2BB2X1 U655 ( .B0(n197), .B1(next_write_addr[6]), .A0N(n198), .A1N(n255), 
        .Y(n259) );
  CLKINVX1 U656 ( .A(write_addr[6]), .Y(n255) );
  OAI221XL U657 ( .A0(n198), .A1(n258), .B0(n257), .B1(n246), .C0(n260), .Y(
        read_addr[5]) );
  CLKINVX1 U658 ( .A(write_addr[5]), .Y(n258) );
  OAI221XL U659 ( .A0(n198), .A1(n262), .B0(n263), .B1(n246), .C0(n264), .Y(
        read_addr[4]) );
  CLKINVX1 U660 ( .A(write_addr[4]), .Y(n262) );
  OAI221XL U661 ( .A0(n198), .A1(n265), .B0(n266), .B1(n246), .C0(n267), .Y(
        read_addr[3]) );
  CLKINVX1 U662 ( .A(write_addr[3]), .Y(n265) );
  OAI221XL U663 ( .A0(n198), .A1(n268), .B0(n269), .B1(n246), .C0(n270), .Y(
        read_addr[2]) );
  CLKINVX1 U664 ( .A(write_addr[2]), .Y(n268) );
  OAI221XL U665 ( .A0(n198), .A1(n271), .B0(n272), .B1(n246), .C0(n273), .Y(
        read_addr[1]) );
  AOI2BB2X1 U666 ( .B0(n261), .B1(next_write_addr[0]), .A0N(n274), .A1N(n195), 
        .Y(n273) );
  CLKINVX1 U667 ( .A(write_addr[1]), .Y(n271) );
  OAI221XL U668 ( .A0(n275), .A1(n196), .B0(n195), .B1(n276), .C0(n277), .Y(
        read_addr[19]) );
  CLKINVX1 U669 ( .A(write_addr[17]), .Y(n276) );
  OAI221XL U670 ( .A0(n279), .A1(n196), .B0(n195), .B1(n280), .C0(n281), .Y(
        read_addr[18]) );
  CLKINVX1 U671 ( .A(write_addr[16]), .Y(n280) );
  OAI221XL U672 ( .A0(n282), .A1(n196), .B0(n195), .B1(n283), .C0(n284), .Y(
        read_addr[17]) );
  OAI221XL U673 ( .A0(n285), .A1(n196), .B0(n195), .B1(n286), .C0(n287), .Y(
        read_addr[16]) );
  OAI221XL U674 ( .A0(n198), .A1(n283), .B0(n282), .B1(n246), .C0(n288), .Y(
        read_addr[15]) );
  CLKINVX1 U675 ( .A(write_addr[15]), .Y(n283) );
  OAI221XL U676 ( .A0(n198), .A1(n286), .B0(n285), .B1(n246), .C0(n290), .Y(
        read_addr[14]) );
  CLKINVX1 U677 ( .A(n195), .Y(n289) );
  CLKINVX1 U678 ( .A(n196), .Y(n261) );
  CLKINVX1 U679 ( .A(write_addr[14]), .Y(n286) );
  OAI221XL U680 ( .A0(n291), .A1(n196), .B0(n195), .B1(n292), .C0(n293), .Y(
        read_addr[13]) );
  CLKINVX1 U681 ( .A(next_write_addr[11]), .Y(n291) );
  OAI221XL U682 ( .A0(n294), .A1(n196), .B0(n195), .B1(n295), .C0(n296), .Y(
        read_addr[12]) );
  CLKINVX1 U683 ( .A(next_write_addr[10]), .Y(n294) );
  OAI221XL U684 ( .A0(n245), .A1(n196), .B0(n244), .B1(n195), .C0(n297), .Y(
        read_addr[11]) );
  AOI2BB2X1 U685 ( .B0(n197), .B1(next_write_addr[11]), .A0N(n198), .A1N(n292), 
        .Y(n297) );
  CLKINVX1 U686 ( .A(write_addr[11]), .Y(n292) );
  CLKINVX1 U687 ( .A(write_addr[9]), .Y(n244) );
  CLKINVX1 U688 ( .A(next_write_addr[9]), .Y(n245) );
  OAI221XL U689 ( .A0(n298), .A1(n196), .B0(n195), .B1(n253), .C0(n299), .Y(
        read_addr[10]) );
  AOI2BB2X1 U690 ( .B0(n197), .B1(next_write_addr[10]), .A0N(n198), .A1N(n295), 
        .Y(n299) );
  CLKINVX1 U691 ( .A(write_addr[10]), .Y(n295) );
  CLKINVX1 U692 ( .A(write_addr[8]), .Y(n253) );
  CLKINVX1 U693 ( .A(n301), .Y(n302) );
  NAND3BX1 U694 ( .AN(n303), .B(n304), .C(n242), .Y(n301) );
  CLKINVX1 U695 ( .A(read_cntr[1]), .Y(n242) );
  CLKINVX1 U696 ( .A(next_write_addr[8]), .Y(n298) );
  AOI21X1 U697 ( .A0(read_cntr[1]), .A1(n311), .B0(n303), .Y(n307) );
  NOR2X1 U698 ( .A(n311), .B(read_cntr[1]), .Y(n303) );
  CLKINVX1 U699 ( .A(read_cntr[0]), .Y(n311) );
  CLKINVX1 U700 ( .A(write_addr[0]), .Y(n274) );
  AOI22X1 U701 ( .A0(N728), .A1(n205), .B0(n199), .B1(write_addr[9]), .Y(n313)
         );
  AO22X1 U702 ( .A0(write_cntr[9]), .A1(n201), .B0(N275), .B1(n316), .Y(
        next_write_cntr[9]) );
  OAI2BB1X1 U703 ( .A0N(next_write_cntr[8]), .A1N(n213), .B0(n317), .Y(
        next_write_addr[8]) );
  AOI22X1 U704 ( .A0(N727), .A1(n205), .B0(write_addr[8]), .B1(n199), .Y(n317)
         );
  OAI2BB1X1 U705 ( .A0N(next_write_cntr[7]), .A1N(n213), .B0(n318), .Y(
        next_write_addr[7]) );
  AOI22X1 U706 ( .A0(N726), .A1(n205), .B0(write_addr[7]), .B1(n199), .Y(n318)
         );
  OAI2BB1X1 U707 ( .A0N(next_write_cntr[6]), .A1N(n213), .B0(n319), .Y(
        next_write_addr[6]) );
  AOI22X1 U708 ( .A0(N725), .A1(n205), .B0(write_addr[6]), .B1(n199), .Y(n319)
         );
  CLKINVX1 U709 ( .A(n263), .Y(next_write_addr[4]) );
  AO22X1 U710 ( .A0(write_cntr[4]), .A1(n201), .B0(N270), .B1(n200), .Y(
        next_write_cntr[4]) );
  CLKINVX1 U711 ( .A(n269), .Y(next_write_addr[2]) );
  AO22X1 U712 ( .A0(n201), .A1(write_cntr[19]), .B0(N285), .B1(n200), .Y(
        next_write_cntr[19]) );
  AO22X1 U713 ( .A0(n201), .A1(write_cntr[18]), .B0(N284), .B1(n316), .Y(
        next_write_cntr[18]) );
  CLKINVX1 U714 ( .A(n275), .Y(next_write_addr[17]) );
  AOI22X1 U715 ( .A0(n38), .A1(n213), .B0(n199), .B1(write_addr[17]), .Y(n275)
         );
  AO22X1 U716 ( .A0(n201), .A1(write_cntr[17]), .B0(N283), .B1(n200), .Y(
        next_write_cntr[17]) );
  CLKINVX1 U717 ( .A(n279), .Y(next_write_addr[16]) );
  AOI22X1 U718 ( .A0(next_write_cntr[16]), .A1(n213), .B0(n199), .B1(
        write_addr[16]), .Y(n279) );
  CLKINVX1 U719 ( .A(n282), .Y(next_write_addr[15]) );
  AOI22X1 U720 ( .A0(next_write_cntr[15]), .A1(n213), .B0(n199), .B1(
        write_addr[15]), .Y(n282) );
  CLKINVX1 U721 ( .A(n285), .Y(next_write_addr[14]) );
  AOI22X1 U722 ( .A0(next_write_cntr[14]), .A1(n213), .B0(n199), .B1(
        write_addr[14]), .Y(n285) );
  OAI2BB1X1 U723 ( .A0N(next_write_cntr[13]), .A1N(n213), .B0(n320), .Y(
        next_write_addr[13]) );
  AOI22X1 U724 ( .A0(N732), .A1(n205), .B0(write_addr[13]), .B1(n199), .Y(n320) );
  OAI2BB1X1 U725 ( .A0N(n41), .A1N(n213), .B0(n321), .Y(next_write_addr[12])
         );
  AOI22X1 U726 ( .A0(N731), .A1(n205), .B0(write_addr[12]), .B1(n199), .Y(n321) );
  AO22X1 U727 ( .A0(write_cntr[12]), .A1(n201), .B0(N278), .B1(n316), .Y(
        next_write_cntr[12]) );
  OAI2BB1X1 U728 ( .A0N(next_write_cntr[11]), .A1N(n213), .B0(n322), .Y(
        next_write_addr[11]) );
  AOI22X1 U729 ( .A0(N730), .A1(n205), .B0(write_addr[11]), .B1(n199), .Y(n322) );
  OAI2BB1X1 U730 ( .A0N(next_write_cntr[10]), .A1N(n213), .B0(n323), .Y(
        next_write_addr[10]) );
  AOI22X1 U731 ( .A0(N729), .A1(n205), .B0(write_addr[10]), .B1(n199), .Y(n323) );
  AO22X1 U732 ( .A0(write_cntr[0]), .A1(n201), .B0(N266), .B1(n200), .Y(
        next_write_cntr[0]) );
  AO22X1 U733 ( .A0(read_cntr[9]), .A1(n203), .B0(N233), .B1(n202), .Y(
        next_read_cntr[9]) );
  AO22X1 U734 ( .A0(read_cntr[8]), .A1(n203), .B0(N232), .B1(n202), .Y(
        next_read_cntr[8]) );
  AO22X1 U735 ( .A0(read_cntr[7]), .A1(n203), .B0(N231), .B1(n202), .Y(
        next_read_cntr[7]) );
  AO22X1 U736 ( .A0(read_cntr[6]), .A1(n203), .B0(N230), .B1(n202), .Y(
        next_read_cntr[6]) );
  AO22X1 U737 ( .A0(read_cntr[5]), .A1(n203), .B0(N229), .B1(n202), .Y(
        next_read_cntr[5]) );
  AO22X1 U738 ( .A0(read_cntr[4]), .A1(n203), .B0(N228), .B1(n202), .Y(
        next_read_cntr[4]) );
  AO22X1 U739 ( .A0(read_cntr[3]), .A1(n203), .B0(N227), .B1(n202), .Y(
        next_read_cntr[3]) );
  AO22X1 U740 ( .A0(read_cntr[2]), .A1(n203), .B0(N226), .B1(n202), .Y(
        next_read_cntr[2]) );
  AO22X1 U741 ( .A0(n203), .A1(read_cntr[1]), .B0(N225), .B1(n202), .Y(
        next_read_cntr[1]) );
  AO22X1 U742 ( .A0(read_cntr[19]), .A1(n203), .B0(N243), .B1(n202), .Y(
        next_read_cntr[19]) );
  AO22X1 U743 ( .A0(read_cntr[18]), .A1(n203), .B0(N242), .B1(n202), .Y(
        next_read_cntr[18]) );
  AO22X1 U744 ( .A0(read_cntr[17]), .A1(n203), .B0(N241), .B1(n202), .Y(
        next_read_cntr[17]) );
  AO22X1 U745 ( .A0(read_cntr[16]), .A1(n203), .B0(N240), .B1(n202), .Y(
        next_read_cntr[16]) );
  AO22X1 U746 ( .A0(read_cntr[15]), .A1(n203), .B0(N239), .B1(n202), .Y(
        next_read_cntr[15]) );
  AO22X1 U747 ( .A0(read_cntr[14]), .A1(n203), .B0(N238), .B1(n202), .Y(
        next_read_cntr[14]) );
  AO22X1 U748 ( .A0(read_cntr[13]), .A1(n203), .B0(N237), .B1(n202), .Y(
        next_read_cntr[13]) );
  AO22X1 U749 ( .A0(read_cntr[12]), .A1(n203), .B0(N236), .B1(n202), .Y(
        next_read_cntr[12]) );
  AO22X1 U750 ( .A0(read_cntr[11]), .A1(n203), .B0(N235), .B1(n202), .Y(
        next_read_cntr[11]) );
  AO22X1 U751 ( .A0(read_cntr[10]), .A1(n203), .B0(N234), .B1(n202), .Y(
        next_read_cntr[10]) );
  AO22X1 U752 ( .A0(n203), .A1(read_cntr[0]), .B0(N224), .B1(n202), .Y(
        next_read_cntr[0]) );
  MXI2X1 U753 ( .A(n340), .B(n341), .S0(n378), .Y(next_photo[1]) );
  OA21XL U754 ( .A0(n342), .A1(curr_photo[0]), .B0(n343), .Y(n340) );
  XOR2X1 U755 ( .A(curr_photo[0]), .B(photo_num[0]), .Y(n345) );
  XNOR2X1 U756 ( .A(n378), .B(photo_num[1]), .Y(n344) );
  AND2X1 U757 ( .A(n346), .B(n13), .Y(n343) );
  CLKINVX1 U758 ( .A(n347), .Y(next_glb_cntr[6]) );
  CLKINVX1 U759 ( .A(n348), .Y(next_glb_cntr[5]) );
  CLKINVX1 U760 ( .A(n349), .Y(next_glb_cntr[1]) );
  CLKINVX1 U761 ( .A(n350), .Y(next_glb_cntr[15]) );
  CLKINVX1 U762 ( .A(n351), .Y(next_glb_cntr[0]) );
  AO22X1 U763 ( .A0(cr_read_cntr[8]), .A1(n352), .B0(N359), .B1(n204), .Y(
        next_cr_read_cntr[8]) );
  AO22X1 U764 ( .A0(cr_read_cntr[7]), .A1(n352), .B0(N358), .B1(n204), .Y(
        next_cr_read_cntr[7]) );
  AO22X1 U765 ( .A0(cr_read_cntr[6]), .A1(n352), .B0(N357), .B1(n204), .Y(
        next_cr_read_cntr[6]) );
  AO22X1 U766 ( .A0(cr_read_cntr[5]), .A1(n352), .B0(N356), .B1(n204), .Y(
        next_cr_read_cntr[5]) );
  AO22X1 U767 ( .A0(cr_read_cntr[4]), .A1(n352), .B0(N355), .B1(n204), .Y(
        next_cr_read_cntr[4]) );
  AO22X1 U768 ( .A0(cr_read_cntr[3]), .A1(n352), .B0(N354), .B1(n204), .Y(
        next_cr_read_cntr[3]) );
  AO22X1 U769 ( .A0(cr_read_cntr[2]), .A1(n352), .B0(N353), .B1(n204), .Y(
        next_cr_read_cntr[2]) );
  AO22X1 U770 ( .A0(cr_read_cntr[1]), .A1(n352), .B0(N352), .B1(n204), .Y(
        next_cr_read_cntr[1]) );
  AO22X1 U771 ( .A0(cr_read_cntr[0]), .A1(n352), .B0(N351), .B1(n204), .Y(
        next_cr_read_cntr[0]) );
  AOI32X1 U772 ( .A0(n354), .A1(n324), .A2(n222), .B0(n353), .B1(n205), .Y(
        n330) );
  CLKINVX1 U773 ( .A(n339), .Y(n354) );
  CLKINVX1 U774 ( .A(n355), .Y(n575) );
  CLKINVX1 U775 ( .A(n356), .Y(n576) );
  CLKINVX1 U776 ( .A(n357), .Y(n577) );
  CLKINVX1 U777 ( .A(n358), .Y(n578) );
  OAI211X1 U778 ( .A0(n446), .A1(n208), .B0(n360), .C0(n361), .Y(n601) );
  AOI22X1 U779 ( .A0(N983), .A1(si_sel), .B0(N1003), .B1(n214), .Y(n361) );
  AOI22X1 U780 ( .A0(N801), .A1(n207), .B0(N781), .B1(n206), .Y(n360) );
  OAI211X1 U781 ( .A0(n447), .A1(n208), .B0(n365), .C0(n366), .Y(n602) );
  AOI22X1 U782 ( .A0(N982), .A1(si_sel), .B0(N1002), .B1(n214), .Y(n366) );
  AOI22X1 U783 ( .A0(N800), .A1(n207), .B0(N780), .B1(n206), .Y(n365) );
  OAI211X1 U784 ( .A0(n448), .A1(n208), .B0(n367), .C0(n368), .Y(n603) );
  AOI22X1 U785 ( .A0(N981), .A1(si_sel), .B0(N1001), .B1(n214), .Y(n368) );
  AOI22X1 U786 ( .A0(N799), .A1(n207), .B0(N779), .B1(n206), .Y(n367) );
  OAI211X1 U787 ( .A0(n449), .A1(n208), .B0(n369), .C0(n370), .Y(n604) );
  AOI22X1 U788 ( .A0(N980), .A1(si_sel), .B0(N1000), .B1(n214), .Y(n370) );
  AOI22X1 U789 ( .A0(N798), .A1(n207), .B0(N778), .B1(n206), .Y(n369) );
  OAI211X1 U790 ( .A0(n450), .A1(n208), .B0(n371), .C0(n372), .Y(n605) );
  AOI22X1 U791 ( .A0(N979), .A1(si_sel), .B0(N999), .B1(n214), .Y(n372) );
  AOI22X1 U792 ( .A0(N797), .A1(n207), .B0(N777), .B1(n206), .Y(n371) );
  OAI211X1 U793 ( .A0(n451), .A1(n208), .B0(n373), .C0(n374), .Y(n606) );
  AOI22X1 U794 ( .A0(N978), .A1(si_sel), .B0(N998), .B1(n214), .Y(n374) );
  AOI22X1 U795 ( .A0(N796), .A1(n207), .B0(N776), .B1(n206), .Y(n373) );
  OAI211X1 U796 ( .A0(n452), .A1(n208), .B0(n375), .C0(n376), .Y(n607) );
  AOI22X1 U797 ( .A0(N977), .A1(si_sel), .B0(N997), .B1(n214), .Y(n376) );
  AOI22X1 U798 ( .A0(N795), .A1(n207), .B0(N775), .B1(n206), .Y(n375) );
  OAI211X1 U799 ( .A0(n453), .A1(n208), .B0(n377), .C0(n380), .Y(n608) );
  AOI22X1 U800 ( .A0(N976), .A1(si_sel), .B0(N996), .B1(n214), .Y(n380) );
  AOI22X1 U801 ( .A0(N976), .A1(n207), .B0(N774), .B1(n206), .Y(n377) );
  OAI211X1 U802 ( .A0(n454), .A1(n208), .B0(n381), .C0(n382), .Y(n609) );
  AOI22X1 U803 ( .A0(N975), .A1(si_sel), .B0(N995), .B1(n214), .Y(n382) );
  AOI22X1 U804 ( .A0(N975), .A1(n207), .B0(N773), .B1(n206), .Y(n381) );
  OAI211X1 U805 ( .A0(n420), .A1(n208), .B0(n383), .C0(n384), .Y(n591) );
  AOI22X1 U806 ( .A0(N993), .A1(si_sel), .B0(N1013), .B1(n214), .Y(n384) );
  AOI22X1 U807 ( .A0(N811), .A1(n207), .B0(N791), .B1(n206), .Y(n383) );
  OAI211X1 U808 ( .A0(n437), .A1(n208), .B0(n385), .C0(n386), .Y(n592) );
  AOI22X1 U809 ( .A0(N992), .A1(si_sel), .B0(N1012), .B1(n214), .Y(n386) );
  AOI22X1 U810 ( .A0(N810), .A1(n207), .B0(N790), .B1(n206), .Y(n385) );
  OAI211X1 U811 ( .A0(n438), .A1(n208), .B0(n387), .C0(n388), .Y(n593) );
  AOI22X1 U812 ( .A0(N991), .A1(si_sel), .B0(N1011), .B1(n214), .Y(n388) );
  AOI22X1 U813 ( .A0(N809), .A1(n207), .B0(N789), .B1(n206), .Y(n387) );
  OAI211X1 U814 ( .A0(n439), .A1(n208), .B0(n389), .C0(n390), .Y(n594) );
  AOI22X1 U815 ( .A0(N990), .A1(si_sel), .B0(N1010), .B1(n214), .Y(n390) );
  AOI22X1 U816 ( .A0(N808), .A1(n207), .B0(N788), .B1(n206), .Y(n389) );
  OAI211X1 U817 ( .A0(n440), .A1(n208), .B0(n391), .C0(n392), .Y(n595) );
  AOI22X1 U818 ( .A0(N989), .A1(si_sel), .B0(N1009), .B1(n214), .Y(n392) );
  AOI22X1 U819 ( .A0(N807), .A1(n207), .B0(N787), .B1(n206), .Y(n391) );
  OAI211X1 U820 ( .A0(n441), .A1(n208), .B0(n393), .C0(n394), .Y(n596) );
  AOI22X1 U821 ( .A0(N988), .A1(si_sel), .B0(N1008), .B1(n214), .Y(n394) );
  AOI22X1 U822 ( .A0(N806), .A1(n207), .B0(N786), .B1(n206), .Y(n393) );
  OAI211X1 U823 ( .A0(n442), .A1(n208), .B0(n395), .C0(n396), .Y(n597) );
  AOI22X1 U824 ( .A0(N987), .A1(si_sel), .B0(N1007), .B1(n214), .Y(n396) );
  AOI22X1 U825 ( .A0(N805), .A1(n207), .B0(N785), .B1(n206), .Y(n395) );
  OAI211X1 U826 ( .A0(n443), .A1(n208), .B0(n397), .C0(n398), .Y(n598) );
  AOI22X1 U827 ( .A0(N986), .A1(si_sel), .B0(N1006), .B1(n214), .Y(n398) );
  AOI22X1 U828 ( .A0(N804), .A1(n207), .B0(N784), .B1(n206), .Y(n397) );
  OAI211X1 U829 ( .A0(n444), .A1(n208), .B0(n399), .C0(n400), .Y(n599) );
  AOI22X1 U830 ( .A0(N985), .A1(si_sel), .B0(N1005), .B1(n214), .Y(n400) );
  AOI22X1 U831 ( .A0(N803), .A1(n207), .B0(N783), .B1(n206), .Y(n399) );
  OAI211X1 U832 ( .A0(n445), .A1(n208), .B0(n401), .C0(n402), .Y(n600) );
  AOI22X1 U833 ( .A0(N984), .A1(si_sel), .B0(N1004), .B1(n214), .Y(n402) );
  AOI22X1 U834 ( .A0(N802), .A1(n207), .B0(N782), .B1(n206), .Y(n401) );
  AOI22X1 U835 ( .A0(N974), .A1(si_sel), .B0(N994), .B1(n214), .Y(n404) );
  AOI22X1 U836 ( .A0(N974), .A1(n207), .B0(N772), .B1(n206), .Y(n403) );
  CLKINVX1 U837 ( .A(n231), .Y(n408) );
  CLKINVX1 U838 ( .A(n410), .Y(n409) );
  AOI21X1 U839 ( .A0(n415), .A1(n416), .B0(n212), .Y(expand_sel[3]) );
  NOR2X1 U840 ( .A(n421), .B(n212), .Y(expand_sel[2]) );
  OAI21XL U841 ( .A0(n217), .A1(n417), .B0(n423), .Y(n422) );
  NOR2X1 U842 ( .A(n424), .B(n212), .Y(expand_sel[1]) );
  OAI21XL U843 ( .A0(N390), .A1(n426), .B0(n417), .Y(n425) );
  NOR2X1 U844 ( .A(n427), .B(n212), .Y(expand_sel[0]) );
  CLKINVX1 U845 ( .A(n429), .Y(n419) );
  MXI2X1 U846 ( .A(n430), .B(n431), .S0(n218), .Y(n428) );
  NOR2X1 U847 ( .A(n230), .B(n426), .Y(n431) );
  NOR2X1 U848 ( .A(n217), .B(n216), .Y(n430) );
  OR2X1 U849 ( .A(n455), .B(n454), .Y(n433) );
  AOI31X1 U850 ( .A0(n435), .A1(n436), .A2(n456), .B0(n212), .Y(n612) );
  AOI222XL U851 ( .A0(N649), .A1(n210), .B0(N667), .B1(n211), .C0(N631), .C1(
        n209), .Y(n456) );
  AOI22X1 U852 ( .A0(N577), .A1(n462), .B0(N613), .B1(n463), .Y(n435) );
  AOI31X1 U853 ( .A0(n464), .A1(n465), .A2(n466), .B0(n212), .Y(n613) );
  AOI222XL U854 ( .A0(N648), .A1(n210), .B0(N666), .B1(n211), .C0(N630), .C1(
        n209), .Y(n466) );
  AOI22X1 U855 ( .A0(N576), .A1(n462), .B0(N612), .B1(n463), .Y(n464) );
  AOI31X1 U856 ( .A0(n468), .A1(n469), .A2(n470), .B0(n212), .Y(n614) );
  AOI222XL U857 ( .A0(N647), .A1(n210), .B0(N665), .B1(n211), .C0(N629), .C1(
        n209), .Y(n470) );
  AOI22X1 U858 ( .A0(N575), .A1(n462), .B0(N611), .B1(n463), .Y(n468) );
  AOI31X1 U859 ( .A0(n471), .A1(n472), .A2(n473), .B0(n212), .Y(n615) );
  AOI222XL U860 ( .A0(N646), .A1(n210), .B0(N664), .B1(n211), .C0(N628), .C1(
        n209), .Y(n473) );
  AOI22X1 U861 ( .A0(N574), .A1(n462), .B0(N610), .B1(n463), .Y(n471) );
  AOI31X1 U862 ( .A0(n474), .A1(n475), .A2(n476), .B0(n212), .Y(n616) );
  AOI222XL U863 ( .A0(N645), .A1(n210), .B0(N663), .B1(n211), .C0(N627), .C1(
        n209), .Y(n476) );
  AOI22X1 U864 ( .A0(N573), .A1(n462), .B0(N609), .B1(n463), .Y(n474) );
  AOI31X1 U865 ( .A0(n477), .A1(n478), .A2(n479), .B0(n212), .Y(n617) );
  AOI222XL U866 ( .A0(N644), .A1(n210), .B0(N662), .B1(n211), .C0(N626), .C1(
        n209), .Y(n479) );
  AOI22X1 U867 ( .A0(N572), .A1(n462), .B0(N608), .B1(n463), .Y(n477) );
  AOI31X1 U868 ( .A0(n480), .A1(n481), .A2(n482), .B0(n212), .Y(n618) );
  AOI222XL U869 ( .A0(N571), .A1(n210), .B0(N571), .B1(n211), .C0(N571), .C1(
        n209), .Y(n482) );
  AOI22X1 U870 ( .A0(N571), .A1(n462), .B0(N571), .B1(n463), .Y(n480) );
  AOI31X1 U871 ( .A0(n483), .A1(n484), .A2(n485), .B0(n212), .Y(n619) );
  AOI222XL U872 ( .A0(N570), .A1(n210), .B0(N570), .B1(n211), .C0(N570), .C1(
        n209), .Y(n485) );
  AOI22X1 U873 ( .A0(N570), .A1(n462), .B0(N570), .B1(n463), .Y(n483) );
  AOI31X1 U874 ( .A0(n486), .A1(n487), .A2(n488), .B0(n212), .Y(n620) );
  AOI222XL U875 ( .A0(N569), .A1(n210), .B0(N569), .B1(n211), .C0(N569), .C1(
        n209), .Y(n488) );
  NOR3X1 U876 ( .A(n211), .B(n210), .C(n209), .Y(n492) );
  AND2X1 U877 ( .A(cr_x[2]), .B(n496), .Y(n493) );
  NAND3X1 U878 ( .A(cr_x[0]), .B(n494), .C(n497), .Y(n489) );
  AOI22X1 U879 ( .A0(N569), .A1(n462), .B0(N569), .B1(n463), .Y(n486) );
  NAND3X1 U880 ( .A(n495), .B(n494), .C(n497), .Y(n490) );
  NOR2BX1 U881 ( .AN(n496), .B(cr_x[2]), .Y(n497) );
  AND2X1 U882 ( .A(n498), .B(n499), .Y(n496) );
  NOR3X1 U883 ( .A(cr_x[6]), .B(cr_x[8]), .C(cr_x[7]), .Y(n499) );
  NOR3X1 U884 ( .A(cr_x[3]), .B(cr_x[5]), .C(cr_x[4]), .Y(n498) );
  CLKINVX1 U885 ( .A(cr_x[0]), .Y(n495) );
  NAND2X1 U886 ( .A(n411), .B(n412), .Y(n405) );
  AOI21X1 U887 ( .A0(N65), .A1(N64), .B0(N66), .Y(n411) );
  NAND2X1 U888 ( .A(n217), .B(n219), .Y(n230) );
  OAI21XL U889 ( .A0(N74), .A1(N73), .B0(N75), .Y(n505) );
  AOI211X1 U890 ( .A0(n507), .A1(n508), .B0(n353), .C0(n237), .Y(n500) );
  AOI211X1 U891 ( .A0(n219), .A1(n216), .B0(n217), .C0(n506), .Y(n237) );
  NOR2X1 U892 ( .A(N76), .B(n429), .Y(n507) );
  NOR4BX1 U893 ( .AN(n509), .B(work_cntr[17]), .C(n74), .D(work_cntr[19]), .Y(
        n429) );
  MXI2X1 U894 ( .A(n512), .B(n513), .S0(n310), .Y(n511) );
  CLKINVX1 U895 ( .A(n412), .Y(n310) );
  NAND2X1 U896 ( .A(curr_photo_size[1]), .B(curr_photo_size[0]), .Y(n412) );
  NAND3BX1 U897 ( .AN(work_cntr[17]), .B(n509), .C(n516), .Y(n506) );
  NOR3X1 U898 ( .A(n74), .B(n218), .C(n85), .Y(n516) );
  AND4X1 U899 ( .A(n517), .B(n518), .C(n519), .D(n520), .Y(n509) );
  NOR4X1 U900 ( .A(n102), .B(n98), .C(n100), .D(n96), .Y(n520) );
  NOR3X1 U901 ( .A(work_cntr[16]), .B(n83), .C(work_cntr[4]), .Y(n519) );
  NOR3X1 U902 ( .A(work_cntr[13]), .B(work_cntr[15]), .C(work_cntr[14]), .Y(
        n518) );
  NOR3X1 U903 ( .A(n76), .B(n92), .C(n88), .Y(n517) );
  CLKINVX1 U904 ( .A(n217), .Y(n306) );
  CLKINVX1 U905 ( .A(n423), .Y(n515) );
  NAND2X1 U906 ( .A(n217), .B(n417), .Y(n423) );
  NAND2X1 U907 ( .A(N390), .B(n426), .Y(n417) );
  CLKINVX1 U908 ( .A(n216), .Y(n426) );
  XOR2X1 U909 ( .A(N82), .B(n521), .Y(n514) );
  NOR2X1 U910 ( .A(N80), .B(N81), .Y(n521) );
  AOI211X1 U911 ( .A0(N87), .A1(N86), .B0(N88), .C0(n522), .Y(n512) );
  NOR3X1 U912 ( .A(N89), .B(N91), .C(N90), .Y(n522) );
  NAND2X1 U913 ( .A(n222), .B(n339), .Y(n329) );
  MXI2X1 U914 ( .A(n523), .B(n524), .S0(si_sel), .Y(n510) );
  CLKINVX1 U915 ( .A(n212), .Y(n621) );
  MXI2X1 U916 ( .A(n527), .B(n528), .S0(N1198), .Y(n524) );
  NAND4BBXL U917 ( .AN(N93), .BN(N92), .C(N95), .D(N94), .Y(n528) );
  NAND4X1 U918 ( .A(n529), .B(n530), .C(n531), .D(n532), .Y(n527) );
  NOR4X1 U919 ( .A(n533), .B(n534), .C(N145), .D(N144), .Y(n532) );
  NAND3X1 U920 ( .A(n331), .B(n337), .C(n332), .Y(n534) );
  CLKINVX1 U921 ( .A(N146), .Y(n332) );
  CLKINVX1 U922 ( .A(N148), .Y(n337) );
  CLKINVX1 U923 ( .A(N147), .Y(n331) );
  CLKINVX1 U924 ( .A(N143), .Y(n333) );
  CLKINVX1 U925 ( .A(N142), .Y(n334) );
  XOR2X1 U926 ( .A(n525), .B(next_state[1]), .Y(n538) );
  MXI2X1 U927 ( .A(n539), .B(n540), .S0(N141), .Y(n535) );
  NAND2X1 U928 ( .A(N139), .B(N140), .Y(n540) );
  NAND2X1 U929 ( .A(n336), .B(n335), .Y(n539) );
  CLKINVX1 U930 ( .A(N140), .Y(n335) );
  CLKINVX1 U931 ( .A(N139), .Y(n336) );
  NOR4X1 U932 ( .A(N152), .B(N151), .C(N150), .D(N149), .Y(n531) );
  NOR3X1 U933 ( .A(N155), .B(N157), .C(N156), .Y(n530) );
  NOR2X1 U934 ( .A(N154), .B(N153), .Y(n529) );
  OAI21XL U935 ( .A0(n13), .A1(n346), .B0(n541), .Y(n523) );
  NOR3X1 U936 ( .A(n573), .B(next_state[1]), .C(n537), .Y(n346) );
  AO21X1 U937 ( .A0(n573), .A1(n537), .B0(n213), .Y(n339) );
  MX3XL U938 ( .A(n13), .B(n547), .C(n544), .S0(n17), .S1(n545), .Y(n546) );
  NAND2X1 U939 ( .A(n548), .B(n526), .Y(n547) );
  MXI2X1 U940 ( .A(n549), .B(n550), .S0(n214), .Y(n548) );
  OAI21XL U941 ( .A0(n551), .A1(n351), .B0(n550), .Y(n549) );
  CLKINVX1 U942 ( .A(n543), .Y(n550) );
  NAND2X1 U943 ( .A(state[2]), .B(n525), .Y(n526) );
  NOR2BX1 U944 ( .AN(n552), .B(n587), .Y(n541) );
  CLKINVX1 U945 ( .A(n551), .Y(n587) );
  NAND2X1 U946 ( .A(N161), .B(n215), .Y(n551) );
  AND3X1 U947 ( .A(n554), .B(n555), .C(n556), .Y(n552) );
  NOR4X1 U948 ( .A(n557), .B(n558), .C(next_glb_cntr[14]), .D(n574), .Y(n556)
         );
  AND2X1 U949 ( .A(N178), .B(n215), .Y(n574) );
  AND2X1 U950 ( .A(N173), .B(n215), .Y(next_glb_cntr[14]) );
  NAND3X1 U951 ( .A(n348), .B(n347), .C(n350), .Y(n558) );
  NAND2X1 U952 ( .A(N174), .B(n215), .Y(n350) );
  NAND2X1 U953 ( .A(N165), .B(n215), .Y(n347) );
  NAND2X1 U954 ( .A(N164), .B(n215), .Y(n348) );
  NAND4X1 U955 ( .A(n358), .B(n357), .C(n356), .D(n355), .Y(n557) );
  NAND2X1 U956 ( .A(N177), .B(n215), .Y(n355) );
  NAND2X1 U957 ( .A(N176), .B(n215), .Y(n356) );
  NAND2X1 U958 ( .A(N175), .B(n215), .Y(n357) );
  NAND2X1 U959 ( .A(N172), .B(n215), .Y(n358) );
  NOR4X1 U960 ( .A(n579), .B(n580), .C(n581), .D(n582), .Y(n555) );
  AND2X1 U961 ( .A(N168), .B(n215), .Y(n582) );
  AND2X1 U962 ( .A(N169), .B(n215), .Y(n581) );
  AND2X1 U963 ( .A(N170), .B(n215), .Y(n580) );
  AND2X1 U964 ( .A(N171), .B(n215), .Y(n579) );
  NOR4X1 U965 ( .A(n583), .B(n584), .C(n585), .D(n586), .Y(n554) );
  AND2X1 U966 ( .A(N162), .B(n215), .Y(n586) );
  AND2X1 U967 ( .A(N163), .B(n215), .Y(n585) );
  AND2X1 U968 ( .A(N166), .B(n215), .Y(n584) );
  AND2X1 U969 ( .A(N167), .B(n215), .Y(n583) );
  NAND2X1 U970 ( .A(N160), .B(n215), .Y(n349) );
  NAND2X1 U971 ( .A(N159), .B(n215), .Y(n351) );
  NOR3X1 U972 ( .A(n446), .B(n451), .C(n450), .Y(n561) );
  NOR3X1 U973 ( .A(n438), .B(n441), .C(n439), .Y(n560) );
  NOR3X1 U974 ( .A(n563), .B(n437), .C(n420), .Y(n559) );
  CLKINVX1 U975 ( .A(n353), .Y(n544) );
  NAND4BX1 U976 ( .AN(write_cntr[12]), .B(n564), .C(n328), .D(n565), .Y(n353)
         );
  OAI31XL U977 ( .A0(n566), .A1(write_cntr[9]), .A2(write_cntr[10]), .B0(
        write_cntr[11]), .Y(n564) );
  CLKINVX1 U978 ( .A(state[2]), .Y(n536) );
  NAND2BX1 U979 ( .AN(n434), .B(n455), .Y(n432) );
  NAND4BX1 U980 ( .AN(n567), .B(n568), .C(n569), .D(n570), .Y(n434) );
  AND2X1 U981 ( .A(n438), .B(n439), .Y(n570) );
  AND3X1 U982 ( .A(n450), .B(n441), .C(n446), .Y(n569) );
  AND2X1 U983 ( .A(n451), .B(n452), .Y(n568) );
  NAND3BX1 U984 ( .AN(n563), .B(n437), .C(n420), .Y(n567) );
  NAND2X1 U985 ( .A(n571), .B(n572), .Y(n563) );
  AND4X1 U986 ( .A(n440), .B(n442), .C(n443), .D(n444), .Y(n572) );
  AND4X1 U987 ( .A(n445), .B(n447), .C(n448), .D(n449), .Y(n571) );
endmodule


module p_dff_WORD24_NSEL5_0 ( clk, reset, en, sel, d, q );
  input [4:0] sel;
  input [23:0] d;
  output [23:0] q;
  input clk, reset, en;
  wire   n50, n51, n76, n77, n78, n79, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n1, n3, n5, n7, n9, n11, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49;

  DFFRHQX1 \q_reg[13]  ( .D(n65), .CK(clk), .RN(n49), .Q(n50) );
  DFFRHQX1 \q_reg[14]  ( .D(n66), .CK(clk), .RN(n49), .Q(q[14]) );
  DFFRHQX1 \q_reg[19]  ( .D(n71), .CK(clk), .RN(n49), .Q(q[19]) );
  DFFRHQX1 \q_reg[17]  ( .D(n69), .CK(clk), .RN(n49), .Q(q[17]) );
  DFFRHQX1 \q_reg[15]  ( .D(n67), .CK(clk), .RN(n49), .Q(q[15]) );
  DFFRHQX1 \q_reg[18]  ( .D(n70), .CK(clk), .RN(n49), .Q(q[18]) );
  DFFRHQX1 \q_reg[16]  ( .D(n68), .CK(clk), .RN(n49), .Q(q[16]) );
  DFFRHQX1 \q_reg[11]  ( .D(n63), .CK(clk), .RN(n49), .Q(n51) );
  DFFRHQX1 \q_reg[3]  ( .D(n55), .CK(clk), .RN(n49), .Q(n78) );
  DFFRHQX1 \q_reg[1]  ( .D(n53), .CK(clk), .RN(n49), .Q(n79) );
  DFFRHQX1 \q_reg[4]  ( .D(n56), .CK(clk), .RN(n49), .Q(n77) );
  DFFRHQX1 \q_reg[10]  ( .D(n62), .CK(clk), .RN(n49), .Q(q[10]) );
  DFFRHQX1 \q_reg[9]  ( .D(n61), .CK(clk), .RN(n49), .Q(n76) );
  DFFRHQX1 \q_reg[2]  ( .D(n54), .CK(clk), .RN(n49), .Q(q[2]) );
  DFFRHQX1 \q_reg[7]  ( .D(n59), .CK(clk), .RN(n49), .Q(q[7]) );
  DFFRHQX1 \q_reg[6]  ( .D(n58), .CK(clk), .RN(n49), .Q(q[6]) );
  DFFRX1 \q_reg[22]  ( .D(n74), .CK(clk), .RN(n49), .Q(q[22]) );
  DFFRX1 \q_reg[21]  ( .D(n73), .CK(clk), .RN(n49), .Q(q[21]) );
  DFFRX1 \q_reg[20]  ( .D(n72), .CK(clk), .RN(n49), .Q(q[20]) );
  DFFRX1 \q_reg[23]  ( .D(n75), .CK(clk), .RN(n49), .Q(q[23]) );
  DFFRHQX2 \q_reg[0]  ( .D(n52), .CK(clk), .RN(n49), .Q(q[0]) );
  DFFRHQX2 \q_reg[5]  ( .D(n57), .CK(clk), .RN(n49), .Q(q[5]) );
  DFFRHQX2 \q_reg[12]  ( .D(n64), .CK(clk), .RN(n49), .Q(q[12]) );
  DFFRHQX2 \q_reg[8]  ( .D(n60), .CK(clk), .RN(n49), .Q(q[8]) );
  MX2XL U3 ( .A(q[16]), .B(d[16]), .S0(n19), .Y(n68) );
  INVXL U4 ( .A(n78), .Y(n1) );
  INVX3 U5 ( .A(n1), .Y(q[3]) );
  INVXL U6 ( .A(n51), .Y(n3) );
  INVX3 U7 ( .A(n3), .Y(q[11]) );
  INVXL U8 ( .A(n50), .Y(n5) );
  INVX3 U9 ( .A(n5), .Y(q[13]) );
  INVXL U10 ( .A(n76), .Y(n7) );
  INVX3 U11 ( .A(n7), .Y(q[9]) );
  INVXL U12 ( .A(n77), .Y(n9) );
  INVX3 U13 ( .A(n9), .Y(q[4]) );
  INVXL U14 ( .A(n79), .Y(n11) );
  INVX3 U15 ( .A(n11), .Y(q[1]) );
  INVX4 U16 ( .A(reset), .Y(n49) );
  OAI21X1 U17 ( .A0(sel[4]), .A1(sel[2]), .B0(n31), .Y(n30) );
  OA21X1 U18 ( .A0(sel[4]), .A1(n22), .B0(n31), .Y(n37) );
  NOR2X2 U19 ( .A(n35), .B(n39), .Y(n31) );
  OAI21X1 U20 ( .A0(sel[3]), .A1(sel[1]), .B0(n16), .Y(n15) );
  OA21X2 U21 ( .A0(sel[3]), .A1(sel[2]), .B0(n19), .Y(n16) );
  INVXL U22 ( .A(n30), .Y(n27) );
  NOR2XL U23 ( .A(n41), .B(n42), .Y(n40) );
  AOI2BB1XL U24 ( .A0N(n22), .A1N(n45), .B0(n35), .Y(n48) );
  AOI2BB1XL U25 ( .A0N(n29), .A1N(sel[1]), .B0(n30), .Y(n28) );
  NOR2XL U26 ( .A(n25), .B(n26), .Y(n24) );
  NOR2XL U27 ( .A(n14), .B(n15), .Y(n13) );
  CLKMX2X2 U28 ( .A(q[23]), .B(d[23]), .S0(n13), .Y(n75) );
  CLKMX2X2 U29 ( .A(d[22]), .B(q[22]), .S0(n15), .Y(n74) );
  CLKMX2X2 U30 ( .A(q[21]), .B(d[21]), .S0(n17), .Y(n73) );
  OA21XL U31 ( .A0(sel[1]), .A1(n18), .B0(n16), .Y(n17) );
  CLKMX2X2 U32 ( .A(q[20]), .B(d[20]), .S0(n16), .Y(n72) );
  CLKMX2X2 U33 ( .A(q[19]), .B(d[19]), .S0(n20), .Y(n71) );
  OA21XL U34 ( .A0(sel[2]), .A1(n18), .B0(n21), .Y(n20) );
  CLKMX2X2 U35 ( .A(q[18]), .B(d[18]), .S0(n21), .Y(n70) );
  OA21XL U36 ( .A0(sel[3]), .A1(n22), .B0(n19), .Y(n21) );
  CLKMX2X2 U37 ( .A(q[17]), .B(d[17]), .S0(n23), .Y(n69) );
  OA21XL U38 ( .A0(n22), .A1(n18), .B0(n19), .Y(n23) );
  CLKINVX1 U39 ( .A(n14), .Y(n18) );
  NOR2X1 U40 ( .A(sel[0]), .B(sel[3]), .Y(n14) );
  AND2X1 U41 ( .A(sel[4]), .B(en), .Y(n19) );
  CLKMX2X2 U42 ( .A(q[15]), .B(d[15]), .S0(n24), .Y(n67) );
  CLKMX2X2 U43 ( .A(d[14]), .B(q[14]), .S0(n26), .Y(n66) );
  OAI21XL U44 ( .A0(sel[4]), .A1(sel[1]), .B0(n27), .Y(n26) );
  CLKMX2X2 U45 ( .A(q[13]), .B(d[13]), .S0(n28), .Y(n65) );
  CLKMX2X2 U46 ( .A(q[12]), .B(d[12]), .S0(n27), .Y(n64) );
  CLKMX2X2 U47 ( .A(q[11]), .B(d[11]), .S0(n32), .Y(n63) );
  AOI21X1 U48 ( .A0(n33), .A1(n34), .B0(n35), .Y(n32) );
  NAND3X1 U49 ( .A(sel[1]), .B(sel[0]), .C(sel[3]), .Y(n34) );
  OAI21XL U50 ( .A0(sel[4]), .A1(sel[2]), .B0(n36), .Y(n33) );
  CLKMX2X2 U51 ( .A(q[10]), .B(d[10]), .S0(n37), .Y(n62) );
  CLKMX2X2 U52 ( .A(q[9]), .B(d[9]), .S0(n38), .Y(n61) );
  OA21XL U53 ( .A0(n22), .A1(n29), .B0(n31), .Y(n38) );
  CLKINVX1 U54 ( .A(n25), .Y(n29) );
  NOR2X1 U55 ( .A(sel[0]), .B(sel[4]), .Y(n25) );
  CLKMX2X2 U56 ( .A(q[8]), .B(d[8]), .S0(n31), .Y(n60) );
  CLKMX2X2 U57 ( .A(q[7]), .B(d[7]), .S0(n40), .Y(n59) );
  CLKMX2X2 U58 ( .A(d[6]), .B(q[6]), .S0(n42), .Y(n58) );
  OAI21XL U59 ( .A0(sel[1]), .A1(n36), .B0(n43), .Y(n42) );
  CLKMX2X2 U60 ( .A(q[5]), .B(d[5]), .S0(n44), .Y(n57) );
  OA21XL U61 ( .A0(sel[1]), .A1(n45), .B0(n43), .Y(n44) );
  CLKMX2X2 U62 ( .A(q[4]), .B(d[4]), .S0(n43), .Y(n56) );
  AOI2BB1X1 U63 ( .A0N(sel[2]), .A1N(n36), .B0(n35), .Y(n43) );
  CLKMX2X2 U64 ( .A(q[3]), .B(d[3]), .S0(n46), .Y(n55) );
  OA21XL U65 ( .A0(sel[2]), .A1(n45), .B0(n47), .Y(n46) );
  CLKMX2X2 U66 ( .A(q[2]), .B(d[2]), .S0(n47), .Y(n54) );
  AOI2BB1X1 U67 ( .A0N(n22), .A1N(n36), .B0(n35), .Y(n47) );
  CLKMX2X2 U68 ( .A(q[1]), .B(d[1]), .S0(n48), .Y(n53) );
  CLKINVX1 U69 ( .A(en), .Y(n35) );
  CLKINVX1 U70 ( .A(n41), .Y(n45) );
  NOR2X1 U71 ( .A(n36), .B(sel[0]), .Y(n41) );
  CLKINVX1 U72 ( .A(n39), .Y(n36) );
  NOR2X1 U73 ( .A(sel[3]), .B(sel[4]), .Y(n39) );
  OR2X1 U74 ( .A(sel[1]), .B(sel[2]), .Y(n22) );
  CLKMX2X2 U75 ( .A(q[0]), .B(d[0]), .S0(en), .Y(n52) );
endmodule


module p_dff_WORD30_NSEL5 ( clk, reset, en, sel, d, q );
  input [4:0] sel;
  input [29:0] d;
  output [29:0] q;
  input clk, reset, en;
  wire   n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n49, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149;

  DFFRXL \q_reg[9]  ( .D(n73), .CK(clk), .RN(n49), .Q(q[9]) );
  DFFRXL \q_reg[19]  ( .D(n83), .CK(clk), .RN(n49), .Q(q[19]) );
  DFFRXL \q_reg[29]  ( .D(n93), .CK(clk), .RN(n49), .Q(q[29]) );
  DFFSRX1 \q_reg[0]  ( .D(n64), .CK(clk), .SN(1'b1), .RN(n149), .QN(n6) );
  DFFSRX1 \q_reg[20]  ( .D(n84), .CK(clk), .SN(1'b1), .RN(n149), .QN(n4) );
  DFFSRX1 \q_reg[10]  ( .D(n74), .CK(clk), .SN(1'b1), .RN(n149), .QN(n5) );
  DFFSRX1 \q_reg[15]  ( .D(n79), .CK(clk), .SN(1'b1), .RN(n149), .QN(n19) );
  DFFSRX1 \q_reg[16]  ( .D(n80), .CK(clk), .SN(1'b1), .RN(n149), .QN(n17) );
  DFFSRX1 \q_reg[17]  ( .D(n81), .CK(clk), .SN(1'b1), .RN(n149), .QN(n18) );
  DFFSRX1 \q_reg[21]  ( .D(n85), .CK(clk), .SN(1'b1), .RN(n149), .QN(n1) );
  DFFSRX1 \q_reg[12]  ( .D(n76), .CK(clk), .SN(1'b1), .RN(n149), .QN(n7) );
  DFFSRX1 \q_reg[11]  ( .D(n75), .CK(clk), .SN(1'b1), .RN(n149), .QN(n3) );
  DFFSRX1 \q_reg[1]  ( .D(n65), .CK(clk), .SN(1'b1), .RN(n149), .QN(n2) );
  DFFSRX1 \q_reg[13]  ( .D(n77), .CK(clk), .SN(1'b1), .RN(n149), .QN(n11) );
  DFFSRX1 \q_reg[26]  ( .D(n90), .CK(clk), .SN(1'b1), .RN(n149), .QN(n22) );
  DFFSRX1 \q_reg[4]  ( .D(n68), .CK(clk), .SN(1'b1), .RN(n149), .QN(n12) );
  DFFSRX1 \q_reg[23]  ( .D(n87), .CK(clk), .SN(1'b1), .RN(n49), .QN(n10) );
  DFFSRX1 \q_reg[24]  ( .D(n88), .CK(clk), .SN(1'b1), .RN(n49), .QN(n14) );
  DFFSRX1 \q_reg[25]  ( .D(n89), .CK(clk), .SN(1'b1), .RN(n49), .QN(n23) );
  DFFSRX1 \q_reg[27]  ( .D(n91), .CK(clk), .SN(1'b1), .RN(n49), .QN(n21) );
  DFFSRX1 \q_reg[2]  ( .D(n66), .CK(clk), .SN(1'b1), .RN(n49), .QN(n8) );
  DFFSRX1 \q_reg[3]  ( .D(n67), .CK(clk), .SN(1'b1), .RN(n49), .QN(n13) );
  DFFSRX1 \q_reg[5]  ( .D(n69), .CK(clk), .SN(1'b1), .RN(n49), .QN(n20) );
  DFFSRX1 \q_reg[7]  ( .D(n71), .CK(clk), .SN(1'b1), .RN(n49), .QN(n16) );
  DFFSRX1 \q_reg[22]  ( .D(n86), .CK(clk), .SN(1'b1), .RN(n149), .QN(n9) );
  DFFSRX1 \q_reg[14]  ( .D(n78), .CK(clk), .SN(1'b1), .RN(n149), .QN(n15) );
  DFFSRX1 \q_reg[6]  ( .D(n70), .CK(clk), .SN(1'b1), .RN(n49), .QN(n24) );
  DFFRX1 \q_reg[8]  ( .D(n72), .CK(clk), .RN(n49), .Q(q[8]) );
  DFFRX1 \q_reg[18]  ( .D(n82), .CK(clk), .RN(n49), .Q(q[18]) );
  DFFRX1 \q_reg[28]  ( .D(n92), .CK(clk), .RN(n49), .Q(q[28]) );
  MX2XL U3 ( .A(q[8]), .B(d[8]), .S0(n131), .Y(n72) );
  INVX16 U4 ( .A(n24), .Y(q[6]) );
  INVX16 U5 ( .A(n15), .Y(q[14]) );
  INVX16 U6 ( .A(n9), .Y(q[22]) );
  INVX16 U7 ( .A(n16), .Y(q[7]) );
  INVX16 U8 ( .A(n20), .Y(q[5]) );
  INVX16 U9 ( .A(n13), .Y(q[3]) );
  INVX16 U10 ( .A(n8), .Y(q[2]) );
  INVX16 U11 ( .A(n21), .Y(q[27]) );
  INVX16 U12 ( .A(n23), .Y(q[25]) );
  INVX16 U13 ( .A(n14), .Y(q[24]) );
  INVX16 U14 ( .A(n10), .Y(q[23]) );
  INVX16 U15 ( .A(n12), .Y(q[4]) );
  INVX16 U16 ( .A(n22), .Y(q[26]) );
  INVX16 U17 ( .A(n11), .Y(q[13]) );
  INVX16 U18 ( .A(n2), .Y(q[1]) );
  INVX16 U19 ( .A(n3), .Y(q[11]) );
  INVX16 U20 ( .A(n7), .Y(q[12]) );
  INVX16 U21 ( .A(n1), .Y(q[21]) );
  INVX16 U22 ( .A(n18), .Y(q[17]) );
  INVX16 U23 ( .A(n17), .Y(q[16]) );
  INVX16 U24 ( .A(n19), .Y(q[15]) );
  INVX16 U25 ( .A(n5), .Y(q[10]) );
  INVX16 U26 ( .A(n4), .Y(q[20]) );
  INVX16 U27 ( .A(n6), .Y(q[0]) );
  CLKBUFX3 U28 ( .A(n149), .Y(n49) );
  INVX3 U29 ( .A(reset), .Y(n149) );
  MX2XL U54 ( .A(q[21]), .B(d[21]), .S0(n118), .Y(n85) );
  MX2XL U55 ( .A(q[1]), .B(d[1]), .S0(n148), .Y(n65) );
  MX2XL U56 ( .A(q[11]), .B(d[11]), .S0(n132), .Y(n75) );
  MX2XL U57 ( .A(d[22]), .B(q[22]), .S0(n116), .Y(n86) );
  MX2XL U58 ( .A(d[6]), .B(q[6]), .S0(n142), .Y(n70) );
  MX2XL U59 ( .A(d[14]), .B(q[14]), .S0(n126), .Y(n78) );
  MX2XL U60 ( .A(q[23]), .B(d[23]), .S0(n114), .Y(n87) );
  MX2XL U61 ( .A(q[7]), .B(d[7]), .S0(n140), .Y(n71) );
  MX2XL U62 ( .A(q[16]), .B(d[16]), .S0(n113), .Y(n80) );
  MX2XL U63 ( .A(q[12]), .B(d[12]), .S0(n127), .Y(n76) );
  MX2XL U64 ( .A(q[2]), .B(d[2]), .S0(n147), .Y(n66) );
  MX2XL U65 ( .A(q[17]), .B(d[17]), .S0(n123), .Y(n81) );
  MX2XL U66 ( .A(q[13]), .B(d[13]), .S0(n128), .Y(n77) );
  MX2XL U67 ( .A(q[15]), .B(d[15]), .S0(n124), .Y(n79) );
  MX2XL U68 ( .A(q[5]), .B(d[5]), .S0(n144), .Y(n69) );
  MX2XL U69 ( .A(q[4]), .B(d[4]), .S0(n143), .Y(n68) );
  MX2XL U70 ( .A(q[27]), .B(d[27]), .S0(n107), .Y(n91) );
  MX2XL U71 ( .A(q[26]), .B(d[26]), .S0(n108), .Y(n90) );
  MX2XL U72 ( .A(q[3]), .B(d[3]), .S0(n146), .Y(n67) );
  MX2XL U73 ( .A(q[25]), .B(d[25]), .S0(n111), .Y(n89) );
  MX2XL U74 ( .A(q[24]), .B(d[24]), .S0(n106), .Y(n88) );
  MX2XL U75 ( .A(q[10]), .B(d[10]), .S0(n137), .Y(n74) );
  MX2XL U76 ( .A(q[20]), .B(d[20]), .S0(n117), .Y(n84) );
  MX2XL U77 ( .A(q[0]), .B(d[0]), .S0(en), .Y(n64) );
  INVX1 U78 ( .A(en), .Y(n135) );
  INVXL U79 ( .A(n130), .Y(n127) );
  CLKMX2X2 U80 ( .A(q[29]), .B(d[29]), .S0(n104), .Y(n93) );
  OA21XL U81 ( .A0(sel[1]), .A1(sel[0]), .B0(n105), .Y(n104) );
  CLKMX2X2 U82 ( .A(q[28]), .B(d[28]), .S0(n105), .Y(n92) );
  AND2X1 U83 ( .A(sel[2]), .B(n106), .Y(n105) );
  OA21XL U84 ( .A0(sel[2]), .A1(sel[0]), .B0(n108), .Y(n107) );
  NOR2X1 U85 ( .A(n109), .B(n110), .Y(n108) );
  AOI2BB1X1 U86 ( .A0N(sel[0]), .A1N(n112), .B0(n109), .Y(n111) );
  CLKINVX1 U87 ( .A(n109), .Y(n106) );
  NAND2X1 U88 ( .A(sel[3]), .B(n113), .Y(n109) );
  NOR2X1 U89 ( .A(n115), .B(n116), .Y(n114) );
  OAI21XL U90 ( .A0(sel[3]), .A1(sel[1]), .B0(n117), .Y(n116) );
  OA21XL U91 ( .A0(sel[1]), .A1(n119), .B0(n117), .Y(n118) );
  AOI2BB1X1 U92 ( .A0N(sel[3]), .A1N(sel[2]), .B0(n120), .Y(n117) );
  CLKMX2X2 U93 ( .A(q[19]), .B(d[19]), .S0(n121), .Y(n83) );
  OA21XL U94 ( .A0(sel[2]), .A1(n119), .B0(n122), .Y(n121) );
  CLKMX2X2 U95 ( .A(q[18]), .B(d[18]), .S0(n122), .Y(n82) );
  AOI2BB1X1 U96 ( .A0N(sel[3]), .A1N(n112), .B0(n120), .Y(n122) );
  AOI2BB1X1 U97 ( .A0N(n119), .A1N(n112), .B0(n120), .Y(n123) );
  CLKINVX1 U98 ( .A(n115), .Y(n119) );
  NOR2X1 U99 ( .A(sel[0]), .B(sel[3]), .Y(n115) );
  CLKINVX1 U100 ( .A(n120), .Y(n113) );
  NAND2X1 U101 ( .A(sel[4]), .B(en), .Y(n120) );
  NOR2X1 U102 ( .A(n125), .B(n126), .Y(n124) );
  OAI21XL U103 ( .A0(sel[4]), .A1(sel[1]), .B0(n127), .Y(n126) );
  AOI2BB1X1 U104 ( .A0N(n129), .A1N(sel[1]), .B0(n130), .Y(n128) );
  OAI21XL U105 ( .A0(sel[4]), .A1(sel[2]), .B0(n131), .Y(n130) );
  AOI21X1 U106 ( .A0(n133), .A1(n134), .B0(n135), .Y(n132) );
  NAND3X1 U107 ( .A(sel[0]), .B(sel[3]), .C(sel[1]), .Y(n134) );
  OAI21XL U108 ( .A0(sel[4]), .A1(sel[2]), .B0(n136), .Y(n133) );
  OA21XL U109 ( .A0(sel[4]), .A1(n112), .B0(n131), .Y(n137) );
  CLKMX2X2 U110 ( .A(q[9]), .B(d[9]), .S0(n138), .Y(n73) );
  OA21XL U111 ( .A0(n112), .A1(n129), .B0(n131), .Y(n138) );
  CLKINVX1 U112 ( .A(n125), .Y(n129) );
  NOR2X1 U113 ( .A(sel[0]), .B(sel[4]), .Y(n125) );
  NOR2X1 U114 ( .A(n135), .B(n139), .Y(n131) );
  NOR2X1 U115 ( .A(n141), .B(n142), .Y(n140) );
  OAI21XL U116 ( .A0(sel[1]), .A1(n136), .B0(n143), .Y(n142) );
  OA21XL U117 ( .A0(sel[1]), .A1(n145), .B0(n143), .Y(n144) );
  AOI2BB1X1 U118 ( .A0N(sel[2]), .A1N(n136), .B0(n135), .Y(n143) );
  OA21XL U119 ( .A0(sel[2]), .A1(n145), .B0(n147), .Y(n146) );
  AOI2BB1X1 U120 ( .A0N(n112), .A1N(n136), .B0(n135), .Y(n147) );
  AOI2BB1X1 U121 ( .A0N(n112), .A1N(n145), .B0(n135), .Y(n148) );
  CLKINVX1 U122 ( .A(n141), .Y(n145) );
  NOR2X1 U123 ( .A(n136), .B(sel[0]), .Y(n141) );
  CLKINVX1 U124 ( .A(n139), .Y(n136) );
  NOR2X1 U125 ( .A(sel[3]), .B(sel[4]), .Y(n139) );
  CLKINVX1 U126 ( .A(n110), .Y(n112) );
  NOR2X1 U127 ( .A(sel[1]), .B(sel[2]), .Y(n110) );
endmodule


module p_dff_WORD24_NSEL5_1 ( clk, reset, en, sel, d, q );
  input [4:0] sel;
  input [23:0] d;
  output [23:0] q;
  input clk, reset, en;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71;

  DFFRX2 \q_reg[18]  ( .D(n43), .CK(clk), .RN(n37), .Q(q[18]) );
  DFFRX2 \q_reg[19]  ( .D(n42), .CK(clk), .RN(n37), .Q(q[19]) );
  DFFRX2 \q_reg[20]  ( .D(n41), .CK(clk), .RN(n37), .Q(q[20]) );
  DFFRX4 \q_reg[21]  ( .D(n40), .CK(clk), .RN(n37), .Q(q[21]) );
  DFFRX4 \q_reg[22]  ( .D(n39), .CK(clk), .RN(n37), .Q(q[22]) );
  DFFRX4 \q_reg[23]  ( .D(n38), .CK(clk), .RN(n37), .Q(q[23]) );
  DFFRX4 \q_reg[13]  ( .D(n48), .CK(clk), .RN(n37), .Q(q[13]) );
  DFFRX4 \q_reg[5]  ( .D(n66), .CK(clk), .RN(n37), .Q(q[5]) );
  DFFRX2 \q_reg[15]  ( .D(n46), .CK(clk), .RN(n37), .Q(q[15]) );
  DFFRX2 \q_reg[14]  ( .D(n47), .CK(clk), .RN(n37), .Q(q[14]) );
  DFFRX2 \q_reg[7]  ( .D(n64), .CK(clk), .RN(n37), .Q(q[7]) );
  DFFRX2 \q_reg[11]  ( .D(n50), .CK(clk), .RN(n37), .Q(q[11]) );
  DFFRX2 \q_reg[6]  ( .D(n65), .CK(clk), .RN(n37), .Q(q[6]) );
  DFFRX2 \q_reg[17]  ( .D(n44), .CK(clk), .RN(n37), .Q(q[17]) );
  DFFRX2 \q_reg[3]  ( .D(n68), .CK(clk), .RN(n37), .Q(q[3]) );
  DFFRX2 \q_reg[10]  ( .D(n51), .CK(clk), .RN(n37), .Q(q[10]) );
  DFFRX2 \q_reg[16]  ( .D(n45), .CK(clk), .RN(n37), .Q(q[16]) );
  DFFRX2 \q_reg[12]  ( .D(n49), .CK(clk), .RN(n37), .Q(q[12]) );
  DFFRX2 \q_reg[9]  ( .D(n62), .CK(clk), .RN(n37), .Q(q[9]) );
  DFFRX2 \q_reg[2]  ( .D(n69), .CK(clk), .RN(n37), .Q(q[2]) );
  DFFRX2 \q_reg[8]  ( .D(n63), .CK(clk), .RN(n37), .Q(q[8]) );
  DFFRX2 \q_reg[4]  ( .D(n67), .CK(clk), .RN(n37), .Q(q[4]) );
  DFFRX2 \q_reg[1]  ( .D(n70), .CK(clk), .RN(n37), .Q(q[1]) );
  DFFRX2 \q_reg[0]  ( .D(n71), .CK(clk), .RN(n37), .Q(q[0]) );
  CLKINVX6 U3 ( .A(reset), .Y(n37) );
  OAI21X1 U4 ( .A0(sel[4]), .A1(sel[2]), .B0(n19), .Y(n18) );
  OA21X1 U5 ( .A0(sel[4]), .A1(n10), .B0(n19), .Y(n25) );
  NOR2X2 U6 ( .A(n23), .B(n27), .Y(n19) );
  OAI21X1 U7 ( .A0(sel[3]), .A1(sel[1]), .B0(n4), .Y(n3) );
  OA21X2 U8 ( .A0(sel[3]), .A1(sel[2]), .B0(n7), .Y(n4) );
  INVX1 U9 ( .A(en), .Y(n23) );
  INVXL U10 ( .A(n18), .Y(n15) );
  NOR2XL U11 ( .A(n29), .B(n30), .Y(n28) );
  AOI2BB1XL U12 ( .A0N(n10), .A1N(n33), .B0(n23), .Y(n36) );
  CLKMX2X2 U13 ( .A(q[23]), .B(d[23]), .S0(n1), .Y(n38) );
  NOR2X1 U14 ( .A(n2), .B(n3), .Y(n1) );
  CLKMX2X2 U15 ( .A(d[22]), .B(q[22]), .S0(n3), .Y(n39) );
  CLKMX2X2 U16 ( .A(q[21]), .B(d[21]), .S0(n5), .Y(n40) );
  OA21XL U17 ( .A0(sel[1]), .A1(n6), .B0(n4), .Y(n5) );
  CLKMX2X2 U18 ( .A(q[20]), .B(d[20]), .S0(n4), .Y(n41) );
  CLKMX2X2 U19 ( .A(q[19]), .B(d[19]), .S0(n8), .Y(n42) );
  OA21XL U20 ( .A0(sel[2]), .A1(n6), .B0(n9), .Y(n8) );
  CLKMX2X2 U21 ( .A(q[18]), .B(d[18]), .S0(n9), .Y(n43) );
  OA21XL U22 ( .A0(sel[3]), .A1(n10), .B0(n7), .Y(n9) );
  CLKMX2X2 U23 ( .A(q[17]), .B(d[17]), .S0(n11), .Y(n44) );
  OA21XL U24 ( .A0(n10), .A1(n6), .B0(n7), .Y(n11) );
  CLKINVX1 U25 ( .A(n2), .Y(n6) );
  NOR2X1 U26 ( .A(sel[0]), .B(sel[3]), .Y(n2) );
  CLKMX2X2 U27 ( .A(q[16]), .B(d[16]), .S0(n7), .Y(n45) );
  AND2X1 U28 ( .A(sel[4]), .B(en), .Y(n7) );
  CLKMX2X2 U29 ( .A(q[15]), .B(d[15]), .S0(n12), .Y(n46) );
  NOR2X1 U30 ( .A(n13), .B(n14), .Y(n12) );
  CLKMX2X2 U31 ( .A(d[14]), .B(q[14]), .S0(n14), .Y(n47) );
  OAI21XL U32 ( .A0(sel[4]), .A1(sel[1]), .B0(n15), .Y(n14) );
  CLKMX2X2 U33 ( .A(q[13]), .B(d[13]), .S0(n16), .Y(n48) );
  AOI2BB1X1 U34 ( .A0N(n17), .A1N(sel[1]), .B0(n18), .Y(n16) );
  CLKMX2X2 U35 ( .A(q[12]), .B(d[12]), .S0(n15), .Y(n49) );
  CLKMX2X2 U36 ( .A(q[11]), .B(d[11]), .S0(n20), .Y(n50) );
  AOI21X1 U37 ( .A0(n21), .A1(n22), .B0(n23), .Y(n20) );
  NAND3X1 U38 ( .A(sel[1]), .B(sel[0]), .C(sel[3]), .Y(n22) );
  OAI21XL U39 ( .A0(sel[4]), .A1(sel[2]), .B0(n24), .Y(n21) );
  CLKMX2X2 U40 ( .A(q[10]), .B(d[10]), .S0(n25), .Y(n51) );
  CLKMX2X2 U41 ( .A(q[9]), .B(d[9]), .S0(n26), .Y(n62) );
  OA21XL U42 ( .A0(n10), .A1(n17), .B0(n19), .Y(n26) );
  CLKINVX1 U43 ( .A(n13), .Y(n17) );
  NOR2X1 U44 ( .A(sel[0]), .B(sel[4]), .Y(n13) );
  CLKMX2X2 U45 ( .A(q[8]), .B(d[8]), .S0(n19), .Y(n63) );
  CLKMX2X2 U46 ( .A(q[7]), .B(d[7]), .S0(n28), .Y(n64) );
  CLKMX2X2 U47 ( .A(d[6]), .B(q[6]), .S0(n30), .Y(n65) );
  OAI21XL U48 ( .A0(sel[1]), .A1(n24), .B0(n31), .Y(n30) );
  CLKMX2X2 U49 ( .A(q[5]), .B(d[5]), .S0(n32), .Y(n66) );
  OA21XL U50 ( .A0(sel[1]), .A1(n33), .B0(n31), .Y(n32) );
  CLKMX2X2 U51 ( .A(q[4]), .B(d[4]), .S0(n31), .Y(n67) );
  AOI2BB1X1 U52 ( .A0N(sel[2]), .A1N(n24), .B0(n23), .Y(n31) );
  CLKMX2X2 U53 ( .A(q[3]), .B(d[3]), .S0(n34), .Y(n68) );
  OA21XL U54 ( .A0(sel[2]), .A1(n33), .B0(n35), .Y(n34) );
  CLKMX2X2 U55 ( .A(q[2]), .B(d[2]), .S0(n35), .Y(n69) );
  AOI2BB1X1 U56 ( .A0N(n10), .A1N(n24), .B0(n23), .Y(n35) );
  CLKMX2X2 U57 ( .A(q[1]), .B(d[1]), .S0(n36), .Y(n70) );
  CLKINVX1 U58 ( .A(n29), .Y(n33) );
  NOR2X1 U59 ( .A(n24), .B(sel[0]), .Y(n29) );
  CLKINVX1 U60 ( .A(n27), .Y(n24) );
  NOR2X1 U61 ( .A(sel[3]), .B(sel[4]), .Y(n27) );
  OR2X1 U62 ( .A(sel[1]), .B(sel[2]), .Y(n10) );
  CLKMX2X2 U63 ( .A(q[0]), .B(d[0]), .S0(en), .Y(n71) );
endmodule


module p_dff_WORD20_NSEL5_2 ( clk, reset, en, sel, d, q );
  input [4:0] sel;
  input [19:0] d;
  output [19:0] q;
  input clk, reset, en;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n52,
         n53, n54, n55, n56, n57, n58, n59;

  DFFRX1 \q_reg[19]  ( .D(n32), .CK(clk), .RN(n31), .Q(q[19]) );
  DFFRX1 \q_reg[0]  ( .D(n59), .CK(clk), .RN(n31), .Q(q[0]) );
  DFFRX1 \q_reg[1]  ( .D(n58), .CK(clk), .RN(n31), .Q(q[1]) );
  DFFRX1 \q_reg[4]  ( .D(n55), .CK(clk), .RN(n31), .Q(q[4]) );
  DFFRX1 \q_reg[2]  ( .D(n57), .CK(clk), .RN(n31), .Q(q[2]) );
  DFFRX1 \q_reg[5]  ( .D(n54), .CK(clk), .RN(n31), .Q(q[5]) );
  DFFRX1 \q_reg[11]  ( .D(n40), .CK(clk), .RN(n31), .Q(q[11]) );
  DFFRX1 \q_reg[6]  ( .D(n53), .CK(clk), .RN(n31), .Q(q[6]) );
  DFFRX1 \q_reg[3]  ( .D(n56), .CK(clk), .RN(n31), .Q(q[3]) );
  DFFRX1 \q_reg[7]  ( .D(n52), .CK(clk), .RN(n31), .Q(q[7]) );
  DFFRX1 \q_reg[16]  ( .D(n35), .CK(clk), .RN(n31), .Q(q[16]) );
  DFFRX1 \q_reg[17]  ( .D(n34), .CK(clk), .RN(n31), .Q(q[17]) );
  DFFRX1 \q_reg[8]  ( .D(n43), .CK(clk), .RN(n31), .Q(q[8]) );
  DFFRX1 \q_reg[10]  ( .D(n41), .CK(clk), .RN(n31), .Q(q[10]) );
  DFFRX1 \q_reg[9]  ( .D(n42), .CK(clk), .RN(n31), .Q(q[9]) );
  DFFRX1 \q_reg[18]  ( .D(n33), .CK(clk), .RN(n31), .Q(q[18]) );
  DFFRX1 \q_reg[12]  ( .D(n39), .CK(clk), .RN(n31), .Q(q[12]) );
  DFFRX1 \q_reg[13]  ( .D(n38), .CK(clk), .RN(n31), .Q(q[13]) );
  DFFRX1 \q_reg[14]  ( .D(n37), .CK(clk), .RN(n31), .Q(q[14]) );
  DFFRX1 \q_reg[15]  ( .D(n36), .CK(clk), .RN(n31), .Q(q[15]) );
  MX2XL U3 ( .A(q[16]), .B(d[16]), .S0(n4), .Y(n35) );
  INVX4 U4 ( .A(reset), .Y(n31) );
  OA21X2 U5 ( .A0(sel[2]), .A1(n18), .B0(en), .Y(n25) );
  INVX1 U6 ( .A(en), .Y(n6) );
  INVXL U7 ( .A(n13), .Y(n10) );
  MX2XL U8 ( .A(d[14]), .B(q[14]), .S0(n9), .Y(n37) );
  MX2XL U9 ( .A(d[12]), .B(q[12]), .S0(n13), .Y(n39) );
  MX2XL U10 ( .A(q[4]), .B(d[4]), .S0(n25), .Y(n55) );
  MX2XL U11 ( .A(q[8]), .B(d[8]), .S0(n14), .Y(n43) );
  MX2XL U12 ( .A(d[6]), .B(q[6]), .S0(n24), .Y(n53) );
  CLKMX2X2 U13 ( .A(d[19]), .B(q[19]), .S0(n1), .Y(n32) );
  OAI31XL U14 ( .A0(sel[2]), .A1(sel[3]), .A2(sel[0]), .B0(n2), .Y(n1) );
  CLKMX2X2 U15 ( .A(q[18]), .B(d[18]), .S0(n2), .Y(n33) );
  OA21XL U16 ( .A0(sel[3]), .A1(n3), .B0(n4), .Y(n2) );
  CLKMX2X2 U17 ( .A(d[17]), .B(q[17]), .S0(n5), .Y(n34) );
  OAI31XL U18 ( .A0(sel[0]), .A1(sel[3]), .A2(n3), .B0(n4), .Y(n5) );
  NOR2BX1 U19 ( .AN(sel[4]), .B(n6), .Y(n4) );
  CLKMX2X2 U20 ( .A(q[15]), .B(d[15]), .S0(n7), .Y(n36) );
  NOR2X1 U21 ( .A(n8), .B(n9), .Y(n7) );
  OAI21XL U22 ( .A0(sel[4]), .A1(sel[1]), .B0(n10), .Y(n9) );
  CLKMX2X2 U23 ( .A(q[13]), .B(d[13]), .S0(n11), .Y(n38) );
  OA21XL U24 ( .A0(n12), .A1(sel[1]), .B0(n10), .Y(n11) );
  OAI21XL U25 ( .A0(sel[4]), .A1(sel[2]), .B0(n14), .Y(n13) );
  CLKMX2X2 U26 ( .A(q[11]), .B(d[11]), .S0(n15), .Y(n40) );
  AOI21X1 U27 ( .A0(n16), .A1(n17), .B0(n6), .Y(n15) );
  NAND3X1 U28 ( .A(sel[1]), .B(sel[0]), .C(sel[3]), .Y(n17) );
  OAI21XL U29 ( .A0(sel[4]), .A1(sel[2]), .B0(n18), .Y(n16) );
  CLKMX2X2 U30 ( .A(q[10]), .B(d[10]), .S0(n19), .Y(n41) );
  OA21XL U31 ( .A0(sel[4]), .A1(n3), .B0(n14), .Y(n19) );
  CLKMX2X2 U32 ( .A(q[9]), .B(d[9]), .S0(n20), .Y(n42) );
  OA21XL U33 ( .A0(n3), .A1(n12), .B0(n14), .Y(n20) );
  CLKINVX1 U34 ( .A(n8), .Y(n12) );
  NOR2X1 U35 ( .A(sel[0]), .B(sel[4]), .Y(n8) );
  NOR2X1 U36 ( .A(n6), .B(n21), .Y(n14) );
  CLKMX2X2 U37 ( .A(q[7]), .B(d[7]), .S0(n22), .Y(n52) );
  NOR2X1 U38 ( .A(n23), .B(n24), .Y(n22) );
  OAI21XL U39 ( .A0(sel[1]), .A1(n18), .B0(n25), .Y(n24) );
  CLKMX2X2 U40 ( .A(q[5]), .B(d[5]), .S0(n26), .Y(n54) );
  OA21XL U41 ( .A0(sel[1]), .A1(n27), .B0(n25), .Y(n26) );
  CLKMX2X2 U42 ( .A(q[3]), .B(d[3]), .S0(n28), .Y(n56) );
  OA21XL U43 ( .A0(sel[2]), .A1(n27), .B0(n29), .Y(n28) );
  CLKMX2X2 U44 ( .A(q[2]), .B(d[2]), .S0(n29), .Y(n57) );
  OA21XL U45 ( .A0(n3), .A1(n18), .B0(en), .Y(n29) );
  CLKMX2X2 U46 ( .A(q[1]), .B(d[1]), .S0(n30), .Y(n58) );
  OA21XL U47 ( .A0(n3), .A1(n27), .B0(en), .Y(n30) );
  CLKINVX1 U48 ( .A(n23), .Y(n27) );
  NOR2X1 U49 ( .A(n18), .B(sel[0]), .Y(n23) );
  CLKINVX1 U50 ( .A(n21), .Y(n18) );
  NOR2X1 U51 ( .A(sel[3]), .B(sel[4]), .Y(n21) );
  OR2X1 U52 ( .A(sel[1]), .B(sel[2]), .Y(n3) );
  CLKMX2X2 U53 ( .A(d[0]), .B(q[0]), .S0(n6), .Y(n59) );
endmodule


module p_dff_WORD2_NSEL5_0 ( clk, reset, en, sel, d, q );
  input [4:0] sel;
  input [1:0] d;
  output [1:0] q;
  input clk, reset, en;
  wire   n5, n6, n7, n8, n2, n3, n4;

  DFFSRX1 \q_reg[0]  ( .D(n7), .CK(clk), .SN(1'b1), .RN(n4), .Q(q[0]), .QN(n2)
         );
  DFFRX1 \q_reg[1]  ( .D(n8), .CK(clk), .RN(n4), .Q(q[1]) );
  CLKINVX1 U3 ( .A(reset), .Y(n4) );
  AO22X1 U4 ( .A0(d[1]), .A1(n3), .B0(q[1]), .B1(n5), .Y(n8) );
  CLKINVX1 U5 ( .A(n5), .Y(n3) );
  OAI31X1 U6 ( .A0(n6), .A1(sel[1]), .A2(sel[0]), .B0(en), .Y(n5) );
  OAI2BB2XL U7 ( .B0(n2), .B1(en), .A0N(d[0]), .A1N(en), .Y(n7) );
  OR3X2 U8 ( .A(sel[4]), .B(sel[3]), .C(sel[2]), .Y(n6) );
endmodule


module p_dff_WORD20_NSEL5_1 ( clk, reset, en, sel, d, q );
  input [4:0] sel;
  input [19:0] d;
  output [19:0] q;
  input clk, reset, en;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n52,
         n53, n54, n55, n56, n57, n58, n59;

  DFFRX1 \q_reg[19]  ( .D(n32), .CK(clk), .RN(n31), .Q(q[19]) );
  DFFRX1 \q_reg[13]  ( .D(n38), .CK(clk), .RN(n31), .Q(q[13]) );
  DFFRX1 \q_reg[10]  ( .D(n41), .CK(clk), .RN(n31), .Q(q[10]) );
  DFFRX1 \q_reg[7]  ( .D(n52), .CK(clk), .RN(n31), .Q(q[7]) );
  DFFRX1 \q_reg[0]  ( .D(n59), .CK(clk), .RN(n31), .Q(q[0]) );
  DFFRX1 \q_reg[1]  ( .D(n58), .CK(clk), .RN(n31), .Q(q[1]) );
  DFFRX1 \q_reg[4]  ( .D(n55), .CK(clk), .RN(n31), .Q(q[4]) );
  DFFRX1 \q_reg[2]  ( .D(n57), .CK(clk), .RN(n31), .Q(q[2]) );
  DFFRX1 \q_reg[5]  ( .D(n54), .CK(clk), .RN(n31), .Q(q[5]) );
  DFFRX1 \q_reg[11]  ( .D(n40), .CK(clk), .RN(n31), .Q(q[11]) );
  DFFRX1 \q_reg[6]  ( .D(n53), .CK(clk), .RN(n31), .Q(q[6]) );
  DFFRX1 \q_reg[3]  ( .D(n56), .CK(clk), .RN(n31), .Q(q[3]) );
  DFFRX1 \q_reg[16]  ( .D(n35), .CK(clk), .RN(n31), .Q(q[16]) );
  DFFRX1 \q_reg[17]  ( .D(n34), .CK(clk), .RN(n31), .Q(q[17]) );
  DFFRX1 \q_reg[8]  ( .D(n43), .CK(clk), .RN(n31), .Q(q[8]) );
  DFFRX1 \q_reg[9]  ( .D(n42), .CK(clk), .RN(n31), .Q(q[9]) );
  DFFRX1 \q_reg[18]  ( .D(n33), .CK(clk), .RN(n31), .Q(q[18]) );
  DFFRX1 \q_reg[12]  ( .D(n39), .CK(clk), .RN(n31), .Q(q[12]) );
  DFFRX1 \q_reg[14]  ( .D(n37), .CK(clk), .RN(n31), .Q(q[14]) );
  DFFRX1 \q_reg[15]  ( .D(n36), .CK(clk), .RN(n31), .Q(q[15]) );
  MX2XL U3 ( .A(q[16]), .B(d[16]), .S0(n4), .Y(n35) );
  INVX4 U4 ( .A(reset), .Y(n31) );
  OA21X2 U5 ( .A0(sel[2]), .A1(n18), .B0(en), .Y(n25) );
  INVX1 U6 ( .A(en), .Y(n6) );
  INVXL U7 ( .A(n13), .Y(n10) );
  MX2XL U8 ( .A(d[14]), .B(q[14]), .S0(n9), .Y(n37) );
  MX2XL U9 ( .A(d[12]), .B(q[12]), .S0(n13), .Y(n39) );
  MX2XL U10 ( .A(q[4]), .B(d[4]), .S0(n25), .Y(n55) );
  MX2XL U11 ( .A(q[8]), .B(d[8]), .S0(n14), .Y(n43) );
  MX2XL U12 ( .A(d[6]), .B(q[6]), .S0(n24), .Y(n53) );
  CLKMX2X2 U13 ( .A(d[19]), .B(q[19]), .S0(n1), .Y(n32) );
  OAI31XL U14 ( .A0(sel[2]), .A1(sel[3]), .A2(sel[0]), .B0(n2), .Y(n1) );
  CLKMX2X2 U15 ( .A(q[18]), .B(d[18]), .S0(n2), .Y(n33) );
  OA21XL U16 ( .A0(sel[3]), .A1(n3), .B0(n4), .Y(n2) );
  CLKMX2X2 U17 ( .A(d[17]), .B(q[17]), .S0(n5), .Y(n34) );
  OAI31XL U18 ( .A0(sel[0]), .A1(sel[3]), .A2(n3), .B0(n4), .Y(n5) );
  NOR2BX1 U19 ( .AN(sel[4]), .B(n6), .Y(n4) );
  CLKMX2X2 U20 ( .A(q[15]), .B(d[15]), .S0(n7), .Y(n36) );
  NOR2X1 U21 ( .A(n8), .B(n9), .Y(n7) );
  OAI21XL U22 ( .A0(sel[4]), .A1(sel[1]), .B0(n10), .Y(n9) );
  CLKMX2X2 U23 ( .A(q[13]), .B(d[13]), .S0(n11), .Y(n38) );
  OA21XL U24 ( .A0(n12), .A1(sel[1]), .B0(n10), .Y(n11) );
  OAI21XL U25 ( .A0(sel[4]), .A1(sel[2]), .B0(n14), .Y(n13) );
  CLKMX2X2 U26 ( .A(q[11]), .B(d[11]), .S0(n15), .Y(n40) );
  AOI21X1 U27 ( .A0(n16), .A1(n17), .B0(n6), .Y(n15) );
  NAND3X1 U28 ( .A(sel[1]), .B(sel[0]), .C(sel[3]), .Y(n17) );
  OAI21XL U29 ( .A0(sel[4]), .A1(sel[2]), .B0(n18), .Y(n16) );
  CLKMX2X2 U30 ( .A(q[10]), .B(d[10]), .S0(n19), .Y(n41) );
  OA21XL U31 ( .A0(sel[4]), .A1(n3), .B0(n14), .Y(n19) );
  CLKMX2X2 U32 ( .A(q[9]), .B(d[9]), .S0(n20), .Y(n42) );
  OA21XL U33 ( .A0(n3), .A1(n12), .B0(n14), .Y(n20) );
  CLKINVX1 U34 ( .A(n8), .Y(n12) );
  NOR2X1 U35 ( .A(sel[0]), .B(sel[4]), .Y(n8) );
  NOR2X1 U36 ( .A(n6), .B(n21), .Y(n14) );
  CLKMX2X2 U37 ( .A(q[7]), .B(d[7]), .S0(n22), .Y(n52) );
  NOR2X1 U38 ( .A(n23), .B(n24), .Y(n22) );
  OAI21XL U39 ( .A0(sel[1]), .A1(n18), .B0(n25), .Y(n24) );
  CLKMX2X2 U40 ( .A(q[5]), .B(d[5]), .S0(n26), .Y(n54) );
  OA21XL U41 ( .A0(sel[1]), .A1(n27), .B0(n25), .Y(n26) );
  CLKMX2X2 U42 ( .A(q[3]), .B(d[3]), .S0(n28), .Y(n56) );
  OA21XL U43 ( .A0(sel[2]), .A1(n27), .B0(n29), .Y(n28) );
  CLKMX2X2 U44 ( .A(q[2]), .B(d[2]), .S0(n29), .Y(n57) );
  OA21XL U45 ( .A0(n3), .A1(n18), .B0(en), .Y(n29) );
  CLKMX2X2 U46 ( .A(q[1]), .B(d[1]), .S0(n30), .Y(n58) );
  OA21XL U47 ( .A0(n3), .A1(n27), .B0(en), .Y(n30) );
  CLKINVX1 U48 ( .A(n23), .Y(n27) );
  NOR2X1 U49 ( .A(n18), .B(sel[0]), .Y(n23) );
  CLKINVX1 U50 ( .A(n21), .Y(n18) );
  NOR2X1 U51 ( .A(sel[3]), .B(sel[4]), .Y(n21) );
  OR2X1 U52 ( .A(sel[1]), .B(sel[2]), .Y(n3) );
  CLKMX2X2 U53 ( .A(d[0]), .B(q[0]), .S0(n6), .Y(n59) );
endmodule


module p_dff_WORD2_NSEL5_1 ( clk, reset, en, sel, d, q );
  input [4:0] sel;
  input [1:0] d;
  output [1:0] q;
  input clk, reset, en;
  wire   n1, n2, n3, n4, n8, n9, n10;

  DFFRX1 \q_reg[0]  ( .D(n8), .CK(clk), .RN(n3), .Q(q[0]) );
  DFFRX1 \q_reg[1]  ( .D(n4), .CK(clk), .RN(n3), .Q(q[1]) );
  CLKINVX1 U2 ( .A(reset), .Y(n3) );
  AO22X1 U3 ( .A0(d[0]), .A1(en), .B0(q[0]), .B1(n2), .Y(n8) );
  INVXL U4 ( .A(en), .Y(n2) );
  AO22X1 U5 ( .A0(d[1]), .A1(n1), .B0(q[1]), .B1(n10), .Y(n4) );
  CLKINVX1 U6 ( .A(n10), .Y(n1) );
  OAI31X1 U7 ( .A0(n9), .A1(sel[1]), .A2(sel[0]), .B0(en), .Y(n10) );
  OR3X2 U8 ( .A(sel[4]), .B(sel[3]), .C(sel[2]), .Y(n9) );
endmodule


module DP_DW01_inc_0 ( A, SUM );
  input [24:0] A;
  output [24:0] SUM;

  wire   [24:2] carry;

  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  XOR2X1 U1_1_23 ( .A(A[23]), .B(carry[23]), .Y(SUM[23]) );
  ADDHXL U1_1_22 ( .A(A[22]), .B(carry[22]), .CO(carry[23]), .S(SUM[22]) );
  ADDHXL U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHXL U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADDHXL U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHXL U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  ADDHXL U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHXL U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  ADDHXL U1_1_20 ( .A(A[20]), .B(carry[20]), .CO(carry[21]), .S(SUM[20]) );
  ADDHXL U1_1_18 ( .A(A[18]), .B(carry[18]), .CO(carry[19]), .S(SUM[18]) );
  ADDHXL U1_1_19 ( .A(A[19]), .B(carry[19]), .CO(carry[20]), .S(SUM[19]) );
  ADDHXL U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  ADDHXL U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  ADDHXL U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHXL U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  ADDHXL U1_1_21 ( .A(A[21]), .B(carry[21]), .CO(carry[22]), .S(SUM[21]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module DP_DW01_inc_1 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  ADDHXL U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHXL U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADDHXL U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHXL U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  XOR2X1 U1 ( .A(carry[15]), .B(A[15]), .Y(SUM[15]) );
  CLKINVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module DP_DW01_inc_2 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  XOR2X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .Y(SUM[7]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module DP_DW01_add_0 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [9:1] carry;

  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  AND2XL U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKXOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XNOR2X1 U3 ( .A(B[9]), .B(n2), .Y(SUM[9]) );
  NAND2X1 U4 ( .A(B[8]), .B(carry[8]), .Y(n2) );
  XOR2X1 U5 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
endmodule


module DP_DW01_add_1 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [9:1] carry;

  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XNOR2X1 U3 ( .A(B[9]), .B(n2), .Y(SUM[9]) );
  NAND2X1 U4 ( .A(B[8]), .B(carry[8]), .Y(n2) );
  XOR2X1 U5 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
endmodule


module DP_DW01_add_2 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [9:1] carry;

  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XNOR2X1 U3 ( .A(B[9]), .B(n2), .Y(SUM[9]) );
  NAND2X1 U4 ( .A(B[8]), .B(carry[8]), .Y(n2) );
  XOR2X1 U5 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
endmodule


module DP ( clk, reset, im_q, cr_q, im_d, en_si, en_init_time, en_fb_addr, 
        en_photo_num, en_curr_photo_addr, en_curr_photo_size, en_so, si_sel, 
        init_time_mux_sel, sftr_n, so_mux_sel, expand_sel, curr_time, fb_addr, 
        photo_num, curr_photo_addr, curr_photo_size );
  input [23:0] im_q;
  input [12:0] cr_q;
  output [29:0] im_d;
  input [1:0] sftr_n;
  input [1:0] so_mux_sel;
  input [3:0] expand_sel;
  output [23:0] curr_time;
  output [19:0] fb_addr;
  output [1:0] photo_num;
  output [19:0] curr_photo_addr;
  output [1:0] curr_photo_size;
  input clk, reset, en_si, en_init_time, en_fb_addr, en_photo_num,
         en_curr_photo_addr, en_curr_photo_size, en_so, si_sel,
         init_time_mux_sel;
  wire   \photo_num_w[1] , N46, N52, N54, N55, N56, N57, N58, N59, N60, N61,
         N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83,
         N84, N85, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122,
         N123, N124, N125, \curr_photo_size_sel[0] , n77, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n63, n64, n65, n69, n71, n72, n73,
         n74, n75, n76, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95;
  wire   [23:0] si_mux;
  wire   [23:0] init_time_mux;
  wire   [23:0] si_w;
  wire   [9:0] addr_b;
  wire   [9:0] addr_g;
  wire   [9:0] addr_r;
  wire   [9:0] sftr_b;
  wire   [9:0] sftr_g;
  wire   [9:0] sftr_r;
  wire   [29:0] so_mux;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;

  NOR4BBX4 U165 ( .AN(N46), .BN(n14), .C(N52), .D(n2), .Y(n157) );
  p_dff_WORD24_NSEL5_0 si_reg ( .clk(clk), .reset(reset), .en(en_si), .sel({
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .d(si_mux), .q(si_w) );
  p_dff_WORD30_NSEL5 so_reg ( .clk(clk), .reset(reset), .en(en_so), .sel({1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1}), .d(so_mux), .q(im_d) );
  p_dff_WORD24_NSEL5_1 init_time_reg ( .clk(clk), .reset(reset), .en(
        en_init_time), .sel({1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .d(init_time_mux), 
        .q(curr_time) );
  p_dff_WORD20_NSEL5_2 fb_addr_reg ( .clk(clk), .reset(reset), .en(en_fb_addr), 
        .sel({1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .d(si_w[19:0]), .q(fb_addr) );
  p_dff_WORD2_NSEL5_0 photo_num_reg ( .clk(clk), .reset(reset), .en(
        en_photo_num), .sel({1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .d({
        \photo_num_w[1] , n19}), .q(photo_num) );
  p_dff_WORD20_NSEL5_1 curr_photo_addr_reg ( .clk(clk), .reset(reset), .en(
        en_curr_photo_addr), .sel({1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .d(
        si_w[19:0]), .q(curr_photo_addr) );
  p_dff_WORD2_NSEL5_1 curr_photo_size_reg ( .clk(clk), .reset(reset), .en(
        en_curr_photo_size), .sel({1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .d({n77, 
        \curr_photo_size_sel[0] }), .q(curr_photo_size) );
  DP_DW01_inc_0 add_125 ( .A({1'b0, curr_time}), .SUM({SYNOPSYS_UNCONNECTED__0, 
        N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, 
        N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102}) );
  DP_DW01_inc_1 add_123 ( .A(curr_time[23:8]), .SUM({N85, N84, N83, N82, N81, 
        N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70}) );
  DP_DW01_inc_2 add_121 ( .A({1'b0, curr_time[23:16]}), .SUM({
        SYNOPSYS_UNCONNECTED__1, N61, N60, N59, N58, N57, N56, N55, N54}) );
  DP_DW01_add_0 add_107 ( .A({1'b0, 1'b0, si_w[23:16]}), .B(im_d[29:20]), .CI(
        1'b0), .SUM(addr_r) );
  DP_DW01_add_1 add_106 ( .A({1'b0, 1'b0, si_w[15:8]}), .B(im_d[19:10]), .CI(
        1'b0), .SUM(addr_g) );
  DP_DW01_add_2 add_105 ( .A({1'b0, 1'b0, si_w[7:0]}), .B(im_d[9:0]), .CI(1'b0), .SUM(addr_b) );
  CLKBUFX2 U3 ( .A(si_sel), .Y(n15) );
  INVXL U4 ( .A(si_w[16]), .Y(n49) );
  AOI32XL U6 ( .A0(curr_time[1]), .A1(curr_time[0]), .A2(curr_time[3]), .B0(
        curr_time[2]), .B1(curr_time[3]), .Y(n22) );
  NOR4XL U7 ( .A(n191), .B(si_w[11]), .C(si_w[13]), .D(si_w[12]), .Y(n186) );
  NOR4XL U8 ( .A(n185), .B(si_w[11]), .C(si_w[13]), .D(si_w[12]), .Y(n180) );
  NOR4XL U9 ( .A(n188), .B(si_w[3]), .C(si_w[5]), .D(si_w[4]), .Y(n187) );
  NOR4XL U10 ( .A(n184), .B(si_w[3]), .C(si_w[5]), .D(si_w[4]), .Y(n183) );
  NAND3XL U11 ( .A(curr_time[16]), .B(curr_time[18]), .C(curr_time[17]), .Y(
        n29) );
  AOI32XL U12 ( .A0(curr_time[9]), .A1(curr_time[8]), .A2(curr_time[11]), .B0(
        curr_time[10]), .B1(curr_time[11]), .Y(n25) );
  INVXL U13 ( .A(expand_sel[1]), .Y(n32) );
  INVXL U14 ( .A(expand_sel[0]), .Y(n31) );
  INVXL U15 ( .A(so_mux_sel[1]), .Y(n35) );
  OR2XL U16 ( .A(n34), .B(so_mux_sel[1]), .Y(n1) );
  NOR2X1 U18 ( .A(n35), .B(n34), .Y(n110) );
  NOR2BX1 U19 ( .AN(n14), .B(N46), .Y(n152) );
  MXI2X1 U20 ( .A(addr_b[8]), .B(addr_b[9]), .S0(sftr_n[0]), .Y(n78) );
  MXI2X1 U21 ( .A(addr_g[8]), .B(addr_g[9]), .S0(sftr_n[0]), .Y(n86) );
  MXI2X1 U22 ( .A(addr_r[8]), .B(addr_r[9]), .S0(sftr_n[0]), .Y(n94) );
  MXI2X1 U23 ( .A(addr_b[6]), .B(addr_b[7]), .S0(sftr_n[0]), .Y(n75) );
  MXI2X1 U24 ( .A(addr_g[6]), .B(addr_g[7]), .S0(sftr_n[0]), .Y(n84) );
  MXI2X1 U27 ( .A(addr_r[6]), .B(addr_r[7]), .S0(sftr_n[0]), .Y(n92) );
  MXI2X1 U29 ( .A(addr_b[2]), .B(addr_b[3]), .S0(sftr_n[0]), .Y(n71) );
  MXI2X1 U30 ( .A(addr_r[2]), .B(addr_r[3]), .S0(sftr_n[0]), .Y(n88) );
  MXI2X1 U31 ( .A(addr_b[4]), .B(addr_b[5]), .S0(sftr_n[0]), .Y(n73) );
  MXI2X1 U32 ( .A(addr_g[4]), .B(addr_g[5]), .S0(sftr_n[0]), .Y(n82) );
  MXI2X1 U33 ( .A(addr_r[4]), .B(addr_r[5]), .S0(sftr_n[0]), .Y(n90) );
  CLKINVX1 U34 ( .A(si_w[10]), .Y(n55) );
  CLKINVX1 U35 ( .A(si_w[6]), .Y(n59) );
  CLKINVX1 U36 ( .A(si_w[0]), .Y(n69) );
  NOR4X1 U37 ( .A(n189), .B(si_w[1]), .C(si_w[21]), .D(si_w[20]), .Y(n182) );
  NOR4X1 U38 ( .A(n190), .B(si_w[14]), .C(si_w[16]), .D(si_w[15]), .Y(n181) );
  CLKBUFX3 U39 ( .A(n110), .Y(n10) );
  CLKBUFX3 U40 ( .A(n110), .Y(n11) );
  CLKBUFX3 U41 ( .A(n109), .Y(n13) );
  CLKBUFX3 U42 ( .A(n109), .Y(n12) );
  CLKBUFX3 U43 ( .A(n111), .Y(n8) );
  CLKBUFX3 U44 ( .A(n111), .Y(n9) );
  INVX3 U45 ( .A(si_sel), .Y(n16) );
  INVX3 U46 ( .A(n18), .Y(n17) );
  NOR2X1 U47 ( .A(n32), .B(n31), .Y(n143) );
  NAND2X1 U48 ( .A(n34), .B(n35), .Y(n111) );
  CLKBUFX3 U49 ( .A(n15), .Y(n18) );
  CLKBUFX3 U50 ( .A(init_time_mux_sel), .Y(n14) );
  NAND2X1 U51 ( .A(expand_sel[1]), .B(n31), .Y(n145) );
  NAND2X1 U52 ( .A(expand_sel[0]), .B(n32), .Y(n146) );
  INVXL U53 ( .A(expand_sel[2]), .Y(n33) );
  NOR2X1 U54 ( .A(expand_sel[1]), .B(expand_sel[0]), .Y(n139) );
  CLKBUFX3 U55 ( .A(n112), .Y(n6) );
  CLKBUFX3 U56 ( .A(n112), .Y(n7) );
  CLKINVX1 U57 ( .A(n1), .Y(n109) );
  CLKINVX1 U58 ( .A(so_mux_sel[0]), .Y(n34) );
  CLKBUFX3 U59 ( .A(n152), .Y(n4) );
  CLKBUFX3 U60 ( .A(n152), .Y(n5) );
  OAI22XL U61 ( .A0(n145), .A1(n55), .B0(n146), .B1(n54), .Y(n149) );
  NAND4XL U62 ( .A(so_mux_sel[1]), .B(n137), .C(n138), .D(n34), .Y(n112) );
  NAND3BXL U63 ( .AN(n139), .B(expand_sel[2]), .C(expand_sel[3]), .Y(n138) );
  OAI2BB2XL U64 ( .B0(n140), .B1(expand_sel[3]), .A0N(expand_sel[3]), .A1N(
        n141), .Y(n137) );
  AOI22X1 U65 ( .A0(N55), .A1(n157), .B0(N119), .B1(n5), .Y(n169) );
  AOI22XL U66 ( .A0(N57), .A1(n157), .B0(N121), .B1(n4), .Y(n165) );
  AOI22XL U67 ( .A0(N59), .A1(n157), .B0(N123), .B1(n4), .Y(n161) );
  CLKINVX1 U68 ( .A(n71), .Y(n37) );
  CLKINVX1 U69 ( .A(n88), .Y(n41) );
  BUFX4 U70 ( .A(n153), .Y(n3) );
  AND3XL U71 ( .A(n2), .B(n14), .C(N46), .Y(n153) );
  OAI22XL U72 ( .A0(n69), .A1(n33), .B0(expand_sel[2]), .B1(n142), .Y(n141) );
  AOI221XL U73 ( .A0(si_w[1]), .A1(n143), .B0(si_w[4]), .B1(n139), .C0(n144), 
        .Y(n142) );
  OAI22XL U74 ( .A0(n145), .A1(n64), .B0(n146), .B1(n63), .Y(n144) );
  OAI211X1 U75 ( .A0(n69), .A1(n8), .B0(n6), .C0(n136), .Y(so_mux[0]) );
  AOI22X1 U76 ( .A0(sftr_b[0]), .A1(n10), .B0(addr_b[0]), .B1(n12), .Y(n136)
         );
  MX3XL U77 ( .A(addr_b[0]), .B(addr_b[1]), .C(n37), .S0(sftr_n[0]), .S1(
        sftr_n[1]), .Y(sftr_b[0]) );
  OAI211X1 U78 ( .A0(n59), .A1(n9), .B0(n7), .C0(n114), .Y(so_mux[6]) );
  AOI22X1 U79 ( .A0(sftr_b[6]), .A1(n10), .B0(addr_b[6]), .B1(n12), .Y(n114)
         );
  MXI2X1 U80 ( .A(n75), .B(n78), .S0(sftr_n[1]), .Y(sftr_b[6]) );
  OAI211X1 U81 ( .A0(n53), .A1(n9), .B0(n6), .C0(n131), .Y(so_mux[14]) );
  AOI22X1 U82 ( .A0(sftr_g[4]), .A1(n11), .B0(addr_g[4]), .B1(n13), .Y(n131)
         );
  MXI2X1 U83 ( .A(n82), .B(n84), .S0(sftr_n[1]), .Y(sftr_g[4]) );
  OAI211X1 U84 ( .A0(n8), .A1(n47), .B0(n6), .C0(n124), .Y(so_mux[22]) );
  AOI22X1 U85 ( .A0(sftr_r[2]), .A1(n10), .B0(addr_r[2]), .B1(n12), .Y(n124)
         );
  MXI2X1 U86 ( .A(n88), .B(n90), .S0(sftr_n[1]), .Y(sftr_r[2]) );
  OAI211X1 U87 ( .A0(n65), .A1(n9), .B0(n6), .C0(n127), .Y(so_mux[1]) );
  AOI22X1 U88 ( .A0(sftr_b[1]), .A1(n11), .B0(addr_b[1]), .B1(n13), .Y(n127)
         );
  OAI211X1 U89 ( .A0(n64), .A1(n9), .B0(n7), .C0(n118), .Y(so_mux[2]) );
  AOI22X1 U90 ( .A0(sftr_b[2]), .A1(n10), .B0(addr_b[2]), .B1(n12), .Y(n118)
         );
  MXI2X1 U91 ( .A(n71), .B(n73), .S0(sftr_n[1]), .Y(sftr_b[2]) );
  OAI211X1 U92 ( .A0(n63), .A1(n9), .B0(n7), .C0(n117), .Y(so_mux[3]) );
  AOI22X1 U93 ( .A0(sftr_b[3]), .A1(n11), .B0(addr_b[3]), .B1(n13), .Y(n117)
         );
  OAI211X1 U94 ( .A0(n61), .A1(n8), .B0(n7), .C0(n116), .Y(so_mux[4]) );
  AOI22X1 U95 ( .A0(sftr_b[4]), .A1(n10), .B0(addr_b[4]), .B1(n12), .Y(n116)
         );
  MXI2X1 U96 ( .A(n73), .B(n75), .S0(sftr_n[1]), .Y(sftr_b[4]) );
  OAI211X1 U97 ( .A0(n60), .A1(n9), .B0(n7), .C0(n115), .Y(so_mux[5]) );
  AOI22X1 U98 ( .A0(sftr_b[5]), .A1(n10), .B0(addr_b[5]), .B1(n12), .Y(n115)
         );
  OAI211X1 U99 ( .A0(n58), .A1(n9), .B0(n7), .C0(n113), .Y(so_mux[7]) );
  AOI22X1 U100 ( .A0(sftr_b[7]), .A1(n10), .B0(addr_b[7]), .B1(n12), .Y(n113)
         );
  OAI211X1 U101 ( .A0(n56), .A1(n9), .B0(n6), .C0(n134), .Y(so_mux[11]) );
  OAI211X1 U102 ( .A0(n55), .A1(n9), .B0(n6), .C0(n133), .Y(so_mux[12]) );
  AOI22X1 U103 ( .A0(sftr_g[2]), .A1(n11), .B0(addr_g[2]), .B1(n13), .Y(n133)
         );
  MXI2X1 U104 ( .A(n80), .B(n82), .S0(sftr_n[1]), .Y(sftr_g[2]) );
  OAI211X1 U105 ( .A0(n54), .A1(n9), .B0(n6), .C0(n132), .Y(so_mux[13]) );
  AOI22X1 U106 ( .A0(sftr_g[3]), .A1(n11), .B0(addr_g[3]), .B1(n13), .Y(n132)
         );
  OAI211X1 U107 ( .A0(n8), .A1(n52), .B0(n6), .C0(n130), .Y(so_mux[15]) );
  AOI22X1 U108 ( .A0(sftr_g[5]), .A1(n11), .B0(addr_g[5]), .B1(n13), .Y(n130)
         );
  OAI211X1 U109 ( .A0(n8), .A1(n51), .B0(n6), .C0(n129), .Y(so_mux[16]) );
  AOI22X1 U110 ( .A0(sftr_g[6]), .A1(n11), .B0(addr_g[6]), .B1(n13), .Y(n129)
         );
  MXI2X1 U111 ( .A(n84), .B(n86), .S0(sftr_n[1]), .Y(sftr_g[6]) );
  OAI211X1 U112 ( .A0(n8), .A1(n50), .B0(n6), .C0(n128), .Y(so_mux[17]) );
  AOI22X1 U113 ( .A0(sftr_g[7]), .A1(n11), .B0(addr_g[7]), .B1(n13), .Y(n128)
         );
  OAI211X1 U114 ( .A0(n8), .A1(n48), .B0(n6), .C0(n125), .Y(so_mux[21]) );
  AOI22X1 U115 ( .A0(sftr_r[1]), .A1(n10), .B0(addr_r[1]), .B1(n13), .Y(n125)
         );
  OAI211X1 U116 ( .A0(n8), .A1(n46), .B0(n7), .C0(n123), .Y(so_mux[23]) );
  AOI22X1 U117 ( .A0(sftr_r[3]), .A1(n10), .B0(addr_r[3]), .B1(n12), .Y(n123)
         );
  OAI211X1 U118 ( .A0(n8), .A1(n45), .B0(n7), .C0(n122), .Y(so_mux[24]) );
  AOI22X1 U119 ( .A0(sftr_r[4]), .A1(n10), .B0(addr_r[4]), .B1(n12), .Y(n122)
         );
  MXI2X1 U120 ( .A(n90), .B(n92), .S0(sftr_n[1]), .Y(sftr_r[4]) );
  OAI211X1 U121 ( .A0(n8), .A1(n44), .B0(n7), .C0(n121), .Y(so_mux[25]) );
  AOI22X1 U122 ( .A0(sftr_r[5]), .A1(n10), .B0(addr_r[5]), .B1(n12), .Y(n121)
         );
  OAI211X1 U123 ( .A0(n8), .A1(n43), .B0(n7), .C0(n120), .Y(so_mux[26]) );
  AOI22X1 U124 ( .A0(sftr_r[6]), .A1(n10), .B0(addr_r[6]), .B1(n12), .Y(n120)
         );
  MXI2X1 U125 ( .A(n92), .B(n94), .S0(sftr_n[1]), .Y(sftr_r[6]) );
  OAI211X1 U126 ( .A0(n8), .A1(n42), .B0(n7), .C0(n119), .Y(so_mux[27]) );
  AOI22X1 U127 ( .A0(sftr_r[7]), .A1(n10), .B0(addr_r[7]), .B1(n12), .Y(n119)
         );
  OAI211X1 U128 ( .A0(n57), .A1(n9), .B0(n6), .C0(n135), .Y(so_mux[10]) );
  AOI22X1 U129 ( .A0(sftr_g[0]), .A1(n11), .B0(addr_g[0]), .B1(n13), .Y(n135)
         );
  OAI211X1 U130 ( .A0(n8), .A1(n49), .B0(n6), .C0(n126), .Y(so_mux[20]) );
  AOI22X1 U131 ( .A0(sftr_r[0]), .A1(n11), .B0(addr_r[0]), .B1(n13), .Y(n126)
         );
  MX3XL U132 ( .A(addr_r[0]), .B(addr_r[1]), .C(n41), .S0(sftr_n[0]), .S1(
        sftr_n[1]), .Y(sftr_r[0]) );
  OA22XL U133 ( .A0(n147), .A1(n33), .B0(expand_sel[2]), .B1(n148), .Y(n140)
         );
  AOI221XL U134 ( .A0(si_w[5]), .A1(n143), .B0(si_w[8]), .B1(n139), .C0(n150), 
        .Y(n147) );
  AOI221XL U135 ( .A0(si_w[9]), .A1(n143), .B0(si_w[12]), .B1(n139), .C0(n149), 
        .Y(n148) );
  OAI22XL U136 ( .A0(n145), .A1(n59), .B0(n146), .B1(n58), .Y(n150) );
  AOI22X1 U137 ( .A0(sftr_g[1]), .A1(n11), .B0(addr_g[1]), .B1(n13), .Y(n134)
         );
  MX3XL U138 ( .A(addr_g[1]), .B(addr_g[2]), .C(n38), .S0(sftr_n[0]), .S1(
        sftr_n[1]), .Y(sftr_g[1]) );
  CLKINVX1 U139 ( .A(n81), .Y(n38) );
  AO22X1 U140 ( .A0(addr_b[8]), .A1(n12), .B0(sftr_b[8]), .B1(n11), .Y(
        so_mux[8]) );
  NOR2X1 U141 ( .A(sftr_n[1]), .B(n78), .Y(sftr_b[8]) );
  AO22X1 U142 ( .A0(addr_g[8]), .A1(n109), .B0(sftr_g[8]), .B1(n11), .Y(
        so_mux[18]) );
  NOR2X1 U143 ( .A(sftr_n[1]), .B(n86), .Y(sftr_g[8]) );
  AO22X1 U144 ( .A0(addr_b[9]), .A1(n13), .B0(sftr_b[9]), .B1(n10), .Y(
        so_mux[9]) );
  NOR2X1 U145 ( .A(sftr_n[1]), .B(n79), .Y(sftr_b[9]) );
  AO22X1 U146 ( .A0(addr_g[9]), .A1(n109), .B0(sftr_g[9]), .B1(n11), .Y(
        so_mux[19]) );
  NOR2X1 U147 ( .A(sftr_n[1]), .B(n87), .Y(sftr_g[9]) );
  AO22X1 U148 ( .A0(addr_r[9]), .A1(n109), .B0(sftr_r[9]), .B1(n11), .Y(
        so_mux[29]) );
  NOR2X1 U149 ( .A(sftr_n[1]), .B(n95), .Y(sftr_r[9]) );
  AO22X1 U150 ( .A0(addr_r[8]), .A1(n13), .B0(sftr_r[8]), .B1(n110), .Y(
        so_mux[28]) );
  NOR2X1 U151 ( .A(sftr_n[1]), .B(n94), .Y(sftr_r[8]) );
  OAI21XL U152 ( .A0(init_time_mux_sel), .A1(n51), .B0(n173), .Y(
        init_time_mux[14]) );
  AOI22X1 U153 ( .A0(N116), .A1(n4), .B0(N76), .B1(n3), .Y(n173) );
  OAI21XL U154 ( .A0(init_time_mux_sel), .A1(n50), .B0(n172), .Y(
        init_time_mux[15]) );
  AOI22X1 U155 ( .A0(N117), .A1(n4), .B0(N77), .B1(n3), .Y(n172) );
  OAI2BB2XL U156 ( .B0(init_time_mux_sel), .B1(n60), .A0N(N107), .A1N(n5), .Y(
        init_time_mux[5]) );
  MXI2X1 U157 ( .A(n76), .B(n79), .S0(sftr_n[1]), .Y(sftr_b[7]) );
  MXI2X1 U158 ( .A(n85), .B(n87), .S0(sftr_n[1]), .Y(sftr_g[7]) );
  MXI2X1 U159 ( .A(n93), .B(n95), .S0(sftr_n[1]), .Y(sftr_r[7]) );
  NAND2BX1 U160 ( .AN(sftr_n[0]), .B(addr_b[9]), .Y(n79) );
  NAND2BX1 U161 ( .AN(sftr_n[0]), .B(addr_g[9]), .Y(n87) );
  NAND2BX1 U162 ( .AN(sftr_n[0]), .B(addr_r[9]), .Y(n95) );
  OAI21XL U163 ( .A0(init_time_mux_sel), .A1(n57), .B0(n154), .Y(
        init_time_mux[8]) );
  AOI22X1 U164 ( .A0(N110), .A1(n4), .B0(N70), .B1(n3), .Y(n154) );
  OAI211X1 U166 ( .A0(n14), .A1(n43), .B0(n158), .C0(n159), .Y(
        init_time_mux[22]) );
  NAND2X1 U167 ( .A(N84), .B(n3), .Y(n158) );
  AOI22XL U168 ( .A0(N60), .A1(n157), .B0(N124), .B1(n4), .Y(n159) );
  OAI2BB2XL U169 ( .B0(init_time_mux_sel), .B1(n59), .A0N(N108), .A1N(n5), .Y(
        init_time_mux[6]) );
  OAI211X1 U170 ( .A0(n14), .A1(n44), .B0(n160), .C0(n161), .Y(
        init_time_mux[21]) );
  NAND2X1 U171 ( .A(N83), .B(n3), .Y(n160) );
  OAI21XL U172 ( .A0(init_time_mux_sel), .A1(n52), .B0(n174), .Y(
        init_time_mux[13]) );
  AOI22X1 U173 ( .A0(N115), .A1(n4), .B0(N75), .B1(n3), .Y(n174) );
  OAI211X1 U174 ( .A0(n14), .A1(n46), .B0(n164), .C0(n165), .Y(
        init_time_mux[19]) );
  NAND2X1 U175 ( .A(N81), .B(n3), .Y(n164) );
  OAI211X1 U176 ( .A0(n14), .A1(n42), .B0(n155), .C0(n156), .Y(
        init_time_mux[23]) );
  NAND2X1 U177 ( .A(N85), .B(n3), .Y(n155) );
  OAI21XL U178 ( .A0(n14), .A1(n56), .B0(n151), .Y(init_time_mux[9]) );
  AOI22X1 U179 ( .A0(N111), .A1(n4), .B0(N71), .B1(n3), .Y(n151) );
  OAI21XL U180 ( .A0(n14), .A1(n55), .B0(n177), .Y(init_time_mux[10]) );
  AOI22X1 U181 ( .A0(N112), .A1(n4), .B0(N72), .B1(n3), .Y(n177) );
  OAI2BB2XL U182 ( .B0(init_time_mux_sel), .B1(n63), .A0N(N105), .A1N(n5), .Y(
        init_time_mux[3]) );
  OAI21XL U183 ( .A0(n14), .A1(n53), .B0(n175), .Y(init_time_mux[12]) );
  AOI22X1 U184 ( .A0(N114), .A1(n4), .B0(N74), .B1(n3), .Y(n175) );
  OAI2BB2XL U185 ( .B0(init_time_mux_sel), .B1(n58), .A0N(N109), .A1N(n5), .Y(
        init_time_mux[7]) );
  OAI21XL U186 ( .A0(init_time_mux_sel), .A1(n54), .B0(n176), .Y(
        init_time_mux[11]) );
  AOI22X1 U187 ( .A0(N113), .A1(n4), .B0(N73), .B1(n3), .Y(n176) );
  OAI2BB2XL U188 ( .B0(init_time_mux_sel), .B1(n65), .A0N(N103), .A1N(n5), .Y(
        init_time_mux[1]) );
  MXI2X1 U189 ( .A(addr_b[3]), .B(addr_b[4]), .S0(sftr_n[0]), .Y(n72) );
  MXI2X1 U190 ( .A(addr_g[3]), .B(addr_g[4]), .S0(sftr_n[0]), .Y(n81) );
  MXI2X1 U191 ( .A(addr_r[3]), .B(addr_r[4]), .S0(sftr_n[0]), .Y(n89) );
  MXI2X1 U192 ( .A(addr_g[2]), .B(addr_g[3]), .S0(sftr_n[0]), .Y(n80) );
  AOI22XL U193 ( .A0(N61), .A1(n157), .B0(N125), .B1(n4), .Y(n156) );
  MXI2X1 U194 ( .A(addr_b[5]), .B(addr_b[6]), .S0(sftr_n[0]), .Y(n74) );
  MXI2X1 U195 ( .A(addr_b[7]), .B(addr_b[8]), .S0(sftr_n[0]), .Y(n76) );
  MXI2X1 U196 ( .A(addr_g[5]), .B(addr_g[6]), .S0(sftr_n[0]), .Y(n83) );
  MXI2X1 U197 ( .A(addr_g[7]), .B(addr_g[8]), .S0(sftr_n[0]), .Y(n85) );
  MXI2X1 U198 ( .A(addr_r[5]), .B(addr_r[6]), .S0(sftr_n[0]), .Y(n91) );
  MXI2X1 U199 ( .A(addr_r[7]), .B(addr_r[8]), .S0(sftr_n[0]), .Y(n93) );
  MXI2X1 U200 ( .A(n72), .B(n74), .S0(sftr_n[1]), .Y(sftr_b[3]) );
  MXI2X1 U201 ( .A(n74), .B(n76), .S0(sftr_n[1]), .Y(sftr_b[5]) );
  MXI2X1 U202 ( .A(n81), .B(n83), .S0(sftr_n[1]), .Y(sftr_g[3]) );
  MXI2X1 U203 ( .A(n83), .B(n85), .S0(sftr_n[1]), .Y(sftr_g[5]) );
  MXI2X1 U204 ( .A(n89), .B(n91), .S0(sftr_n[1]), .Y(sftr_r[3]) );
  MXI2X1 U205 ( .A(n91), .B(n93), .S0(sftr_n[1]), .Y(sftr_r[5]) );
  OAI211X1 U206 ( .A0(n14), .A1(n45), .B0(n162), .C0(n163), .Y(
        init_time_mux[20]) );
  NAND2X1 U207 ( .A(N82), .B(n3), .Y(n162) );
  AOI22XL U208 ( .A0(N58), .A1(n157), .B0(N122), .B1(n4), .Y(n163) );
  AND2X2 U209 ( .A(im_q[20]), .B(n16), .Y(si_mux[20]) );
  AO22X1 U210 ( .A0(im_q[8]), .A1(n17), .B0(cr_q[8]), .B1(n15), .Y(si_mux[8])
         );
  AND2X2 U211 ( .A(im_q[22]), .B(n16), .Y(si_mux[22]) );
  AO22X1 U212 ( .A0(im_q[6]), .A1(n16), .B0(cr_q[6]), .B1(n15), .Y(si_mux[6])
         );
  AND2X2 U213 ( .A(im_q[14]), .B(n16), .Y(si_mux[14]) );
  OAI2BB2XL U214 ( .B0(init_time_mux_sel), .B1(n61), .A0N(N106), .A1N(n5), .Y(
        init_time_mux[4]) );
  AO22X1 U215 ( .A0(im_q[4]), .A1(n17), .B0(cr_q[4]), .B1(n15), .Y(si_mux[4])
         );
  OAI211X1 U216 ( .A0(n14), .A1(n47), .B0(n166), .C0(n167), .Y(
        init_time_mux[18]) );
  NAND2X1 U217 ( .A(N80), .B(n3), .Y(n166) );
  AOI22XL U218 ( .A0(N56), .A1(n157), .B0(N120), .B1(n5), .Y(n167) );
  AND2X2 U219 ( .A(im_q[18]), .B(n16), .Y(si_mux[18]) );
  OAI211X1 U220 ( .A0(n14), .A1(n49), .B0(n170), .C0(n171), .Y(
        init_time_mux[16]) );
  NAND2X1 U221 ( .A(N78), .B(n3), .Y(n170) );
  AOI22XL U222 ( .A0(N54), .A1(n157), .B0(N118), .B1(n5), .Y(n171) );
  AND2X2 U223 ( .A(im_q[16]), .B(n16), .Y(si_mux[16]) );
  OAI2BB2XL U224 ( .B0(init_time_mux_sel), .B1(n64), .A0N(N104), .A1N(n5), .Y(
        init_time_mux[2]) );
  OAI211X1 U225 ( .A0(n14), .A1(n48), .B0(n168), .C0(n169), .Y(
        init_time_mux[17]) );
  NAND2X1 U226 ( .A(N79), .B(n3), .Y(n168) );
  AO22X1 U227 ( .A0(im_q[9]), .A1(n17), .B0(n18), .B1(cr_q[9]), .Y(si_mux[9])
         );
  AND2X2 U228 ( .A(im_q[21]), .B(n16), .Y(si_mux[21]) );
  AO22X1 U229 ( .A0(im_q[5]), .A1(n17), .B0(cr_q[5]), .B1(n15), .Y(si_mux[5])
         );
  AND2X2 U230 ( .A(im_q[17]), .B(n16), .Y(si_mux[17]) );
  AND2X2 U231 ( .A(im_q[19]), .B(n16), .Y(si_mux[19]) );
  AO22X1 U232 ( .A0(im_q[3]), .A1(n17), .B0(cr_q[3]), .B1(n15), .Y(si_mux[3])
         );
  AND2X2 U233 ( .A(im_q[23]), .B(n16), .Y(si_mux[23]) );
  AND2X2 U234 ( .A(im_q[13]), .B(n16), .Y(si_mux[13]) );
  AO22X1 U235 ( .A0(im_q[7]), .A1(n17), .B0(cr_q[7]), .B1(n15), .Y(si_mux[7])
         );
  AND2X2 U236 ( .A(im_q[15]), .B(n16), .Y(si_mux[15]) );
  AO22X1 U237 ( .A0(im_q[0]), .A1(n16), .B0(cr_q[0]), .B1(n15), .Y(si_mux[0])
         );
  MX3XL U238 ( .A(addr_b[1]), .B(addr_b[2]), .C(n36), .S0(sftr_n[0]), .S1(
        sftr_n[1]), .Y(sftr_b[1]) );
  CLKINVX1 U239 ( .A(n72), .Y(n36) );
  MX3XL U240 ( .A(addr_r[1]), .B(addr_r[2]), .C(n40), .S0(sftr_n[0]), .S1(
        sftr_n[1]), .Y(sftr_r[1]) );
  CLKINVX1 U241 ( .A(n89), .Y(n40) );
  MX3XL U242 ( .A(addr_g[0]), .B(addr_g[1]), .C(n39), .S0(sftr_n[0]), .S1(
        sftr_n[1]), .Y(sftr_g[0]) );
  CLKINVX1 U243 ( .A(n80), .Y(n39) );
  AO22X1 U244 ( .A0(im_q[1]), .A1(n17), .B0(cr_q[1]), .B1(n18), .Y(si_mux[1])
         );
  AO22X1 U245 ( .A0(im_q[2]), .A1(n17), .B0(cr_q[2]), .B1(si_sel), .Y(
        si_mux[2]) );
  AO22X1 U246 ( .A0(im_q[10]), .A1(n17), .B0(cr_q[10]), .B1(n15), .Y(
        si_mux[10]) );
  AO22X1 U247 ( .A0(im_q[11]), .A1(n17), .B0(cr_q[11]), .B1(n15), .Y(
        si_mux[11]) );
  AO22X1 U248 ( .A0(im_q[12]), .A1(n17), .B0(cr_q[12]), .B1(n15), .Y(
        si_mux[12]) );
  CLKINVX1 U249 ( .A(curr_time[21]), .Y(n30) );
  AO22X1 U250 ( .A0(n25), .A1(n24), .B0(n24), .B1(n23), .Y(n2) );
  OAI2BB2XL U251 ( .B0(init_time_mux_sel), .B1(n69), .A0N(N102), .A1N(n5), .Y(
        init_time_mux[0]) );
  NAND2X1 U252 ( .A(n178), .B(n179), .Y(\curr_photo_size_sel[0] ) );
  NAND4X1 U253 ( .A(n180), .B(n181), .C(n182), .D(n183), .Y(n179) );
  CLKINVX1 U254 ( .A(n178), .Y(n77) );
  CLKINVX1 U255 ( .A(si_w[7]), .Y(n58) );
  CLKINVX1 U256 ( .A(si_w[2]), .Y(n64) );
  CLKINVX1 U257 ( .A(si_w[3]), .Y(n63) );
  CLKINVX1 U258 ( .A(si_w[11]), .Y(n54) );
  NAND3X1 U259 ( .A(n42), .B(n64), .C(n43), .Y(n189) );
  NAND3X1 U260 ( .A(n47), .B(n46), .C(n48), .Y(n190) );
  NAND3X1 U261 ( .A(n57), .B(n56), .C(n59), .Y(n184) );
  NAND3X1 U262 ( .A(n69), .B(n55), .C(si_w[7]), .Y(n185) );
  CLKINVX1 U263 ( .A(si_w[8]), .Y(n57) );
  NAND4X1 U264 ( .A(n186), .B(n181), .C(n182), .D(n187), .Y(n178) );
  NAND3X1 U265 ( .A(n58), .B(n57), .C(n59), .Y(n188) );
  CLKINVX1 U266 ( .A(si_w[9]), .Y(n56) );
  CLKINVX1 U267 ( .A(si_w[4]), .Y(n61) );
  CLKINVX1 U268 ( .A(si_w[5]), .Y(n60) );
  CLKINVX1 U269 ( .A(si_w[12]), .Y(n53) );
  CLKINVX1 U270 ( .A(si_w[1]), .Y(n65) );
  CLKINVX1 U271 ( .A(si_w[13]), .Y(n52) );
  CLKINVX1 U272 ( .A(si_w[17]), .Y(n48) );
  CLKINVX1 U273 ( .A(si_w[19]), .Y(n46) );
  CLKINVX1 U274 ( .A(si_w[18]), .Y(n47) );
  CLKINVX1 U275 ( .A(si_w[22]), .Y(n43) );
  CLKINVX1 U276 ( .A(si_w[23]), .Y(n42) );
  CLKINVX1 U277 ( .A(si_w[15]), .Y(n50) );
  CLKINVX1 U278 ( .A(si_w[14]), .Y(n51) );
  NAND3X1 U279 ( .A(n69), .B(n55), .C(si_w[9]), .Y(n191) );
  CLKINVX1 U280 ( .A(si_w[20]), .Y(n45) );
  CLKINVX1 U281 ( .A(si_w[21]), .Y(n44) );
  CLKINVX1 U282 ( .A(si_w[0]), .Y(n19) );
  XOR2X1 U283 ( .A(n19), .B(si_w[1]), .Y(\photo_num_w[1] ) );
  NOR2X1 U284 ( .A(curr_time[7]), .B(curr_time[6]), .Y(n21) );
  NAND2X1 U285 ( .A(curr_time[5]), .B(curr_time[4]), .Y(n20) );
  AOI22X1 U286 ( .A0(n22), .A1(n21), .B0(n21), .B1(n20), .Y(N46) );
  NOR2X1 U287 ( .A(curr_time[15]), .B(curr_time[14]), .Y(n24) );
  NAND2X1 U288 ( .A(curr_time[13]), .B(curr_time[12]), .Y(n23) );
  OR2X1 U289 ( .A(curr_time[23]), .B(curr_time[22]), .Y(n26) );
  NOR2X1 U290 ( .A(curr_time[19]), .B(n26), .Y(n28) );
  NOR3X1 U291 ( .A(n26), .B(curr_time[21]), .C(curr_time[20]), .Y(n27) );
  AOI31X1 U292 ( .A0(n29), .A1(n30), .A2(n28), .B0(n27), .Y(N52) );
endmodule


module DPA ( clk, reset, IM_A, IM_Q, IM_D, IM_WEN, CR_A, CR_Q );
  output [19:0] IM_A;
  input [23:0] IM_Q;
  output [23:0] IM_D;
  output [8:0] CR_A;
  input [12:0] CR_Q;
  input clk, reset;
  output IM_WEN;
  wire   en_si, en_init_time, en_fb_addr, en_photo_num, en_curr_photo_addr,
         en_curr_photo_size, en_so, si_sel, init_time_mux_sel, n1, n2;
  wire   [23:0] curr_time;
  wire   [19:0] fb_addr;
  wire   [1:0] photo_num;
  wire   [19:0] curr_photo_addr;
  wire   [1:0] curr_photo_size;
  wire   [1:0] sftr_n;
  wire   [1:0] so_mux_sel;
  wire   [3:0] expand_sel;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5;

  CONT ctrl_logic ( .clk(clk), .reset(n1), .im_a(IM_A), .im_wen_n(IM_WEN), 
        .cr_a(CR_A), .curr_time(curr_time), .fb_addr(fb_addr), .photo_num(
        photo_num), .curr_photo_addr(curr_photo_addr), .curr_photo_size(
        curr_photo_size), .en_si(en_si), .en_init_time(en_init_time), 
        .en_fb_addr(en_fb_addr), .en_photo_num(en_photo_num), 
        .en_curr_photo_addr(en_curr_photo_addr), .en_curr_photo_size(
        en_curr_photo_size), .en_so(en_so), .si_sel(si_sel), 
        .init_time_mux_sel(init_time_mux_sel), .so_mux_sel(so_mux_sel), 
        .expand_sel(expand_sel) );
  DP data_path ( .clk(clk), .reset(n1), .im_q(IM_Q), .cr_q(CR_Q), .im_d({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, IM_D[23:16], 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, IM_D[15:8], 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, IM_D[7:0]}), .en_si(
        en_si), .en_init_time(en_init_time), .en_fb_addr(en_fb_addr), 
        .en_photo_num(en_photo_num), .en_curr_photo_addr(en_curr_photo_addr), 
        .en_curr_photo_size(en_curr_photo_size), .en_so(en_so), .si_sel(si_sel), .init_time_mux_sel(n2), .sftr_n({1'b1, 1'b0}), .so_mux_sel(so_mux_sel), 
        .expand_sel(expand_sel), .curr_time(curr_time), .fb_addr(fb_addr), 
        .photo_num(photo_num), .curr_photo_addr(curr_photo_addr), 
        .curr_photo_size(curr_photo_size) );
  BUFX4 U1 ( .A(reset), .Y(n1) );
  CLKBUFX3 U2 ( .A(init_time_mux_sel), .Y(n2) );
endmodule

